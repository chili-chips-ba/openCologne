`timescale 1ns / 1ps
module dummy_tb;
    initial begin
        $display("Hello, Verilator!");
        $finish;
    end
endmodule
