mem['h0000] = 32'h00000517;
mem['h0001] = 32'h78050513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'hFF060613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFD050513;
mem['h000E] = 32'h84818593;
mem['h000F] = 32'h00B55863;
mem['h0010] = 32'h00052023;
mem['h0011] = 32'h00450513;
mem['h0012] = 32'hFEB54CE3;
mem['h0013] = 32'h10008117;
mem['h0014] = 32'hFB410113;
mem['h0015] = 32'h10000197;
mem['h0016] = 32'h7AC18193;
mem['h0017] = 32'h00A54533;
mem['h0018] = 32'h00B5C5B3;
mem['h0019] = 32'h00C64633;
mem['h001A] = 32'h6AC000EF;
mem['h001B] = 32'h0000006F;
mem['h001C] = 32'h00000793;
mem['h001D] = 32'h00C79463;
mem['h001E] = 32'h00008067;
mem['h001F] = 32'h00F58733;
mem['h0020] = 32'h00074683;
mem['h0021] = 32'h00F50733;
mem['h0022] = 32'h00178793;
mem['h0023] = 32'h00D70023;
mem['h0024] = 32'hFE5FF06F;
mem['h0025] = 32'h00054783;
mem['h0026] = 32'h0005C703;
mem['h0027] = 32'h00E79463;
mem['h0028] = 32'h00079663;
mem['h0029] = 32'h40E78533;
mem['h002A] = 32'h00008067;
mem['h002B] = 32'h00150513;
mem['h002C] = 32'h00158593;
mem['h002D] = 32'hFE1FF06F;
mem['h002E] = 32'h00251793;
mem['h002F] = 32'h40A78533;
mem['h0030] = 32'h00008067;
mem['h0031] = 32'h200007B7;
mem['h0032] = 32'h0007A703;
mem['h0033] = 32'hFE074EE3;
mem['h0034] = 32'h00A78023;
mem['h0035] = 32'h00008067;
mem['h0036] = 32'hFF010113;
mem['h0037] = 32'h00812423;
mem['h0038] = 32'h01212023;
mem['h0039] = 32'hFFF58413;
mem['h003A] = 32'h00912223;
mem['h003B] = 32'h00112623;
mem['h003C] = 32'h00050493;
mem['h003D] = 32'h00241413;
mem['h003E] = 32'h73C00913;
mem['h003F] = 32'h00045E63;
mem['h0040] = 32'h00C12083;
mem['h0041] = 32'h00812403;
mem['h0042] = 32'h00412483;
mem['h0043] = 32'h00012903;
mem['h0044] = 32'h01010113;
mem['h0045] = 32'h00008067;
mem['h0046] = 32'h0084D7B3;
mem['h0047] = 32'h00F7F793;
mem['h0048] = 32'h00F907B3;
mem['h0049] = 32'h0007C503;
mem['h004A] = 32'hFFC40413;
mem['h004B] = 32'hF99FF0EF;
mem['h004C] = 32'hFCDFF06F;
mem['h004D] = 32'hFF010113;
mem['h004E] = 32'h00812423;
mem['h004F] = 32'h00112623;
mem['h0050] = 32'h00050413;
mem['h0051] = 32'h00044503;
mem['h0052] = 32'h00051A63;
mem['h0053] = 32'h00C12083;
mem['h0054] = 32'h00812403;
mem['h0055] = 32'h01010113;
mem['h0056] = 32'h00008067;
mem['h0057] = 32'h00140413;
mem['h0058] = 32'hF65FF0EF;
mem['h0059] = 32'hFE1FF06F;
mem['h005A] = 32'h20000637;
mem['h005B] = 32'h00462783;
mem['h005C] = 32'h00078F13;
mem['h005D] = 32'h1A07D663;
mem['h005E] = 32'h400006B7;
mem['h005F] = 32'h00D7F6B3;
mem['h0060] = 32'h00068A63;
mem['h0061] = 32'h82018A23;
mem['h0062] = 32'h00100793;
mem['h0063] = 32'h02F60423;
mem['h0064] = 32'h00008067;
mem['h0065] = 32'h0FF7F793;
mem['h0066] = 32'h02400593;
mem['h0067] = 32'h04B79E63;
mem['h0068] = 32'h83418793;
mem['h0069] = 32'h0017C683;
mem['h006A] = 32'h0FF00793;
mem['h006B] = 32'h00F69663;
mem['h006C] = 32'h00200793;
mem['h006D] = 32'hFD9FF06F;
mem['h006E] = 32'h8341C683;
mem['h006F] = 32'h00F69663;
mem['h0070] = 32'h00300793;
mem['h0071] = 32'h02F60423;
mem['h0072] = 32'hFFF00793;
mem['h0073] = 32'h82F18A23;
mem['h0074] = 32'h82018E23;
mem['h0075] = 32'h100007B7;
mem['h0076] = 32'h00078793;
mem['h0077] = 32'h00079023;
mem['h0078] = 32'h0007A223;
mem['h0079] = 32'h0007A423;
mem['h007A] = 32'h0007A623;
mem['h007B] = 32'h200007B7;
mem['h007C] = 32'h02078423;
mem['h007D] = 32'h00008067;
mem['h007E] = 32'h8341C583;
mem['h007F] = 32'h00059663;
mem['h0080] = 32'h00400793;
mem['h0081] = 32'hF89FF06F;
mem['h0082] = 32'h00D00613;
mem['h0083] = 32'h02C78063;
mem['h0084] = 32'h02C00613;
mem['h0085] = 32'h00C78C63;
mem['h0086] = 32'h00A00693;
mem['h0087] = 32'h0CD79063;
mem['h0088] = 32'hF0000793;
mem['h0089] = 32'h82F19A23;
mem['h008A] = 32'h00008067;
mem['h008B] = 32'h100007B7;
mem['h008C] = 32'h00078713;
mem['h008D] = 32'h00174703;
mem['h008E] = 32'h00300613;
mem['h008F] = 32'h00078793;
mem['h0090] = 32'h0EE66063;
mem['h0091] = 32'h83C1CE03;
mem['h0092] = 32'h8201AC23;
mem['h0093] = 32'h00000813;
mem['h0094] = 32'h00000313;
mem['h0095] = 32'h00060513;
mem['h0096] = 32'h84018893;
mem['h0097] = 32'h0FF87613;
mem['h0098] = 32'h03C66E63;
mem['h0099] = 32'h00030463;
mem['h009A] = 32'h82D1AC23;
mem['h009B] = 32'h00200613;
mem['h009C] = 32'h8381A683;
mem['h009D] = 32'h04C70C63;
mem['h009E] = 32'h00300613;
mem['h009F] = 32'h04C70C63;
mem['h00A0] = 32'h00100613;
mem['h00A1] = 32'h04C70063;
mem['h00A2] = 32'h00D78023;
mem['h00A3] = 32'h00170713;
mem['h00A4] = 32'h82018E23;
mem['h00A5] = 32'h00E780A3;
mem['h00A6] = 32'h00008067;
mem['h00A7] = 32'h01180633;
mem['h00A8] = 32'h00064303;
mem['h00A9] = 32'h00269613;
mem['h00AA] = 32'h00D606B3;
mem['h00AB] = 32'h00169693;
mem['h00AC] = 32'hFD068693;
mem['h00AD] = 32'h00D306B3;
mem['h00AE] = 32'h00180813;
mem['h00AF] = 32'h00100313;
mem['h00B0] = 32'hF9DFF06F;
mem['h00B1] = 32'h00D7A223;
mem['h00B2] = 32'hFC5FF06F;
mem['h00B3] = 32'h00D7A423;
mem['h00B4] = 32'hFBDFF06F;
mem['h00B5] = 32'h00D7A623;
mem['h00B6] = 32'hFB5FF06F;
mem['h00B7] = 32'hFD078693;
mem['h00B8] = 32'h0FF6F693;
mem['h00B9] = 32'h00900613;
mem['h00BA] = 32'h00D66863;
mem['h00BB] = 32'h83C1C683;
mem['h00BC] = 32'h00700593;
mem['h00BD] = 32'h00D5FC63;
mem['h00BE] = 32'h82018A23;
mem['h00BF] = 32'h200007B7;
mem['h00C0] = 32'h00500713;
mem['h00C1] = 32'h02E78423;
mem['h00C2] = 32'h00008067;
mem['h00C3] = 32'h00168713;
mem['h00C4] = 32'h82E18E23;
mem['h00C5] = 32'h84018713;
mem['h00C6] = 32'h00D70733;
mem['h00C7] = 32'h00F70023;
mem['h00C8] = 32'h00008067;
mem['h00C9] = 32'h83418793;
mem['h00CA] = 32'h0017C703;
mem['h00CB] = 32'h0C070463;
mem['h00CC] = 32'h000780A3;
mem['h00CD] = 32'h100007B7;
mem['h00CE] = 32'h00078793;
mem['h00CF] = 32'h0017C683;
mem['h00D0] = 32'h00300713;
mem['h00D1] = 32'h00E68A63;
mem['h00D2] = 32'h200007B7;
mem['h00D3] = 32'h00600713;
mem['h00D4] = 32'h02E78423;
mem['h00D5] = 32'h00008067;
mem['h00D6] = 32'h0007C703;
mem['h00D7] = 32'h0ED70863;
mem['h00D8] = 32'h02E6E463;
mem['h00D9] = 32'h00100613;
mem['h00DA] = 32'h02C70E63;
mem['h00DB] = 32'h00200693;
mem['h00DC] = 32'h08D70463;
mem['h00DD] = 32'h00B00713;
mem['h00DE] = 32'h200007B7;
mem['h00DF] = 32'h02E78423;
mem['h00E0] = 32'h00300713;
mem['h00E1] = 32'h06C0006F;
mem['h00E2] = 32'h00400693;
mem['h00E3] = 32'hFED714E3;
mem['h00E4] = 32'h200006B7;
mem['h00E5] = 32'h0246A703;
mem['h00E6] = 32'h10075663;
mem['h00E7] = 32'h00A00793;
mem['h00E8] = 32'h0BC0006F;
mem['h00E9] = 32'h8281C603;
mem['h00EA] = 32'h0FF00713;
mem['h00EB] = 32'h00E61863;
mem['h00EC] = 32'h200007B7;
mem['h00ED] = 32'h00700713;
mem['h00EE] = 32'hF99FF06F;
mem['h00EF] = 32'h0087A703;
mem['h00F0] = 32'h0047A783;
mem['h00F1] = 32'h00F71713;
mem['h00F2] = 32'h01179793;
mem['h00F3] = 32'h0117D793;
mem['h00F4] = 32'h00F767B3;
mem['h00F5] = 32'h82F19823;
mem['h00F6] = 32'h8301A703;
mem['h00F7] = 32'h200007B7;
mem['h00F8] = 32'h00E7A423;
mem['h00F9] = 32'hFFF00713;
mem['h00FA] = 32'h82E18423;
mem['h00FB] = 32'h00200713;
mem['h00FC] = 32'h00E78C23;
mem['h00FD] = 32'h00008067;
mem['h00FE] = 32'h82818693;
mem['h00FF] = 32'h0016C583;
mem['h0100] = 32'h0FF00713;
mem['h0101] = 32'h00E59863;
mem['h0102] = 32'h200007B7;
mem['h0103] = 32'h00800713;
mem['h0104] = 32'hF41FF06F;
mem['h0105] = 32'h0087A703;
mem['h0106] = 32'h0047A783;
mem['h0107] = 32'h00F71713;
mem['h0108] = 32'h01179793;
mem['h0109] = 32'h0117D793;
mem['h010A] = 32'h00F767B3;
mem['h010B] = 32'h82F19823;
mem['h010C] = 32'h8301A703;
mem['h010D] = 32'h200007B7;
mem['h010E] = 32'h00E7A823;
mem['h010F] = 32'hFFF00713;
mem['h0110] = 32'h00E680A3;
mem['h0111] = 32'h00C78C23;
mem['h0112] = 32'h00008067;
mem['h0113] = 32'h200006B7;
mem['h0114] = 32'h0206A703;
mem['h0115] = 32'h00075863;
mem['h0116] = 32'h00900793;
mem['h0117] = 32'h02F68423;
mem['h0118] = 32'h00008067;
mem['h0119] = 32'h0047A703;
mem['h011A] = 32'h0087A783;
mem['h011B] = 32'h03FF05B7;
mem['h011C] = 32'h01071713;
mem['h011D] = 32'h00B77733;
mem['h011E] = 32'h01179793;
mem['h011F] = 32'h82C1A583;
mem['h0120] = 32'h0117D793;
mem['h0121] = 32'h00F767B3;
mem['h0122] = 32'hFC008737;
mem['h0123] = 32'h00B77733;
mem['h0124] = 32'h00E7E7B3;
mem['h0125] = 32'h82F1A623;
mem['h0126] = 32'h02F6A023;
mem['h0127] = 32'h00068C23;
mem['h0128] = 32'h00008067;
mem['h0129] = 32'h0047A703;
mem['h012A] = 32'h0087A783;
mem['h012B] = 32'h03FF05B7;
mem['h012C] = 32'h01071713;
mem['h012D] = 32'h00B77733;
mem['h012E] = 32'h01179793;
mem['h012F] = 32'h82C1A583;
mem['h0130] = 32'h0117D793;
mem['h0131] = 32'h00F767B3;
mem['h0132] = 32'hFC008737;
mem['h0133] = 32'h00B77733;
mem['h0134] = 32'h00E7E7B3;
mem['h0135] = 32'h82F1A623;
mem['h0136] = 32'h02F6A223;
mem['h0137] = 32'hFC1FF06F;
mem['h0138] = 32'h82818693;
mem['h0139] = 32'h0026D603;
mem['h013A] = 32'h82818713;
mem['h013B] = 32'h08061063;
mem['h013C] = 32'h8281C603;
mem['h013D] = 32'h0FF00793;
mem['h013E] = 32'h02F61C63;
mem['h013F] = 32'h200007B7;
mem['h0140] = 32'h0087A603;
mem['h0141] = 32'h02064663;
mem['h0142] = 32'h00C7A703;
mem['h0143] = 32'h82E1A223;
mem['h0144] = 32'h00100713;
mem['h0145] = 32'h82E18023;
mem['h0146] = 32'h40000737;
mem['h0147] = 32'h80E1AC23;
mem['h0148] = 32'h80018E23;
mem['h0149] = 32'hFFF00793;
mem['h014A] = 32'h00F68123;
mem['h014B] = 32'h00008067;
mem['h014C] = 32'h00174683;
mem['h014D] = 32'h0FF00793;
mem['h014E] = 32'h02F69A63;
mem['h014F] = 32'h200007B7;
mem['h0150] = 32'h0107A683;
mem['h0151] = 32'h0206C463;
mem['h0152] = 32'h0147A683;
mem['h0153] = 32'h82D1A223;
mem['h0154] = 32'h00200693;
mem['h0155] = 32'h82D18023;
mem['h0156] = 32'h404006B7;
mem['h0157] = 32'h80D1AC23;
mem['h0158] = 32'h80018E23;
mem['h0159] = 32'hFFF00793;
mem['h015A] = 32'h00F701A3;
mem['h015B] = 32'h00008067;
mem['h015C] = 32'h200007B7;
mem['h015D] = 32'h0007A783;
mem['h015E] = 32'h1807CC63;
mem['h015F] = 32'h82818793;
mem['h0160] = 32'h0027D703;
mem['h0161] = 32'h18070663;
mem['h0162] = 32'hFF010113;
mem['h0163] = 32'h00812423;
mem['h0164] = 32'h81C1C703;
mem['h0165] = 32'h00112623;
mem['h0166] = 32'h00B00613;
mem['h0167] = 32'h02E66E63;
mem['h0168] = 32'h00271713;
mem['h0169] = 32'h75000613;
mem['h016A] = 32'h00C70733;
mem['h016B] = 32'h00072703;
mem['h016C] = 32'h00070067;
mem['h016D] = 32'h200007B7;
mem['h016E] = 32'h02400713;
mem['h016F] = 32'h00E78023;
mem['h0170] = 32'h0180006F;
mem['h0171] = 32'h8201C783;
mem['h0172] = 32'h20000737;
mem['h0173] = 32'h03078793;
mem['h0174] = 32'h0FF7F793;
mem['h0175] = 32'h00F70023;
mem['h0176] = 32'h81C1C783;
mem['h0177] = 32'h00C12083;
mem['h0178] = 32'h00178793;
mem['h0179] = 32'h80F18E23;
mem['h017A] = 32'h00812403;
mem['h017B] = 32'h01010113;
mem['h017C] = 32'h00008067;
mem['h017D] = 32'h200007B7;
mem['h017E] = 32'h02C00713;
mem['h017F] = 32'hFC1FF06F;
mem['h0180] = 32'h8241A503;
mem['h0181] = 32'h00F51513;
mem['h0182] = 32'h00F55513;
mem['h0183] = 32'hAADFF0EF;
mem['h0184] = 32'h82A1A023;
mem['h0185] = 32'h01055513;
mem['h0186] = 32'h00200593;
mem['h0187] = 32'h0FF57513;
mem['h0188] = 32'h00C0006F;
mem['h0189] = 32'h8211C503;
mem['h018A] = 32'h00200593;
mem['h018B] = 32'hAADFF0EF;
mem['h018C] = 32'hFA9FF06F;
mem['h018D] = 32'h8201C503;
mem['h018E] = 32'h00200593;
mem['h018F] = 32'hFF1FF06F;
mem['h0190] = 32'h200007B7;
mem['h0191] = 32'h02C00713;
mem['h0192] = 32'h00E78023;
mem['h0193] = 32'h8001A823;
mem['h0194] = 32'hF89FF06F;
mem['h0195] = 32'h8181A783;
mem['h0196] = 32'h0007A503;
mem['h0197] = 32'h80A1AA23;
mem['h0198] = 32'hFB5FF06F;
mem['h0199] = 32'h8151C503;
mem['h019A] = 32'h00200593;
mem['h019B] = 32'hFC1FF06F;
mem['h019C] = 32'h8141C503;
mem['h019D] = 32'h00200593;
mem['h019E] = 32'hA61FF0EF;
mem['h019F] = 32'h8101A703;
mem['h01A0] = 32'h00170713;
mem['h01A1] = 32'h80E1A823;
mem['h01A2] = 32'h8181A783;
mem['h01A3] = 32'h00478793;
mem['h01A4] = 32'h80F1AC23;
mem['h01A5] = 32'h8241A783;
mem['h01A6] = 32'h00F79793;
mem['h01A7] = 32'h00F7D793;
mem['h01A8] = 32'hF2F70CE3;
mem['h01A9] = 32'h00600793;
mem['h01AA] = 32'h80F18E23;
mem['h01AB] = 32'hF2DFF06F;
mem['h01AC] = 32'h20000737;
mem['h01AD] = 32'h00D00613;
mem['h01AE] = 32'h00C70023;
mem['h01AF] = 32'h0027C603;
mem['h01B0] = 32'h0FF00713;
mem['h01B1] = 32'h00E61463;
mem['h01B2] = 32'h82018423;
mem['h01B3] = 32'h0037C683;
mem['h01B4] = 32'h0FF00713;
mem['h01B5] = 32'hF0E692E3;
mem['h01B6] = 32'h000780A3;
mem['h01B7] = 32'hEFDFF06F;
mem['h01B8] = 32'h20000737;
mem['h01B9] = 32'h00A00693;
mem['h01BA] = 32'h00D70023;
mem['h01BB] = 32'h0027C683;
mem['h01BC] = 32'h0FF00713;
mem['h01BD] = 32'h00E69463;
mem['h01BE] = 32'h00078123;
mem['h01BF] = 32'h0037C683;
mem['h01C0] = 32'h0FF00713;
mem['h01C1] = 32'hECE69AE3;
mem['h01C2] = 32'h000781A3;
mem['h01C3] = 32'hECDFF06F;
mem['h01C4] = 32'h00008067;
mem['h01C5] = 32'hFF010113;
mem['h01C6] = 32'h00112623;
mem['h01C7] = 32'h200007B7;
mem['h01C8] = 32'h00300713;
mem['h01C9] = 32'h00E78C23;
mem['h01CA] = 32'hA41FF0EF;
mem['h01CB] = 32'hBF9FF0EF;
mem['h01CC] = 32'hDB1FF0EF;
mem['h01CD] = 32'hE3DFF0EF;
mem['h01CE] = 32'hFF1FF06F;
mem['h01CF] = 32'h33323130;
mem['h01D0] = 32'h37363534;
mem['h01D1] = 32'h42413938;
mem['h01D2] = 32'h46454443;
mem['h01D3] = 32'h00000000;
mem['h01D4] = 32'h000005B4;
mem['h01D5] = 32'h000005C4;
mem['h01D6] = 32'h000005F4;
mem['h01D7] = 32'h00000600;
mem['h01D8] = 32'h00000624;
mem['h01D9] = 32'h00000634;
mem['h01DA] = 32'h00000640;
mem['h01DB] = 32'h00000654;
mem['h01DC] = 32'h00000664;
mem['h01DD] = 32'h00000670;
mem['h01DE] = 32'h000006B0;
mem['h01DF] = 32'h000006E0;
