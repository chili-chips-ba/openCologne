//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 July 2024)
//  Compile Time: 2024-07-19 13:57:40
//  Program Run:  2024-08-25 18:25:00
//  Program Call: /home/user/FPGA/Boards/GateMate/cc-toolchain-linux//bin/p_r/p_r -i net/top_checkered_synth.v -o top_checkered -ccf top_checkered.ccf -cCP 
//  File Type:    Verilog

// Gatecount:   1076
module top_checkered (btn , clk ,
       led , oled_clk , oled_clk_1 , oled_csn , oled_dc , oled_dc_1 , 
       oled_mosi , oled_mosi_1 , oled_resn , oled_resn_1 
       ) ;

input  btn;
input  clk;

output led;
output oled_clk;
output oled_clk_1;
output oled_csn;
output oled_dc;
output oled_dc_1;
output oled_mosi;
output oled_mosi_1;
output oled_resn;
output oled_resn_1;



wire btn;
wire clk;
wire led;
wire na1_2;
wire na6_1;
wire na7_1;
wire na8_2;
wire na10_1;
wire na11_1;
wire na11_2;
wire na12_1;
wire na13_1;
wire na13_2;
wire na14_1;
wire na17_1;
wire na17_2;
wire na19_1;
wire na19_2;
wire na20_2;
wire na21_1;
wire na22_1;
wire na23_1;
wire na25_1;
wire na29_1;
wire na30_1;
wire na31_1;
wire na32_1;
wire na35_1;
wire na36_1;
wire na39_2;
wire na44_1;
wire na48_1;
wire na48_2;
wire na49_1;
wire na51_1;
wire na51_1_i;
wire na51_2;
wire na51_2_i;
wire na54_1;
wire na55_1;
wire na56_1;
wire na57_2;
wire na58_1;
wire na61_1;
wire na62_1;
wire na63_1;
wire na63_1_i;
wire na63_2;
wire na63_2_i;
wire na64_1;
wire na66_1;
wire na66_1_i;
wire na69_2;
wire na70_1;
wire na72_1;
wire na73_1;
wire na74_2;
wire na74_2_i;
wire na75_1;
wire na77_1;
wire na78_1;
wire na78_1_i;
wire na78_2;
wire na78_2_i;
wire na79_1;
wire na80_1;
wire na80_1_i;
wire na80_2;
wire na80_2_i;
wire na81_1;
wire na83_2;
wire na83_2_i;
wire na84_1;
wire na85_1;
wire na87_1;
wire na88_1;
wire na89_1;
wire na89_1_i;
wire na89_2;
wire na89_2_i;
wire na90_1;
wire na92_2;
wire na92_2_i;
wire na93_1;
wire na94_1;
wire na95_1;
wire na95_1_i;
wire na96_1;
wire na96_2;
wire na97_1;
wire na98_2;
wire na99_2;
wire na99_2_i;
wire na100_1;
wire na102_1;
wire na102_1_i;
wire na103_1;
wire na104_1;
wire na106_1;
wire na107_2;
wire na109_1;
wire na110_1;
wire na111_2;
wire na111_2_i;
wire na112_1;
wire na115_1;
wire na117_1;
wire na117_1_i;
wire na118_1;
wire na119_1;
wire na121_2;
wire na121_2_i;
wire na122_1;
wire na123_1;
wire na125_2;
wire na127_1;
wire na128_1;
wire na130_1;
wire na131_1;
wire na131_1_i;
wire na131_2;
wire na131_2_i;
wire na132_1;
wire na133_1;
wire na133_1_i;
wire na134_1;
wire na135_1;
wire na135_1_i;
wire na135_2;
wire na135_2_i;
wire na136_2;
wire na137_1;
wire na137_2;
wire na138_1;
wire na138_2;
wire na139_1;
wire na139_2;
wire na141_1;
wire na141_2;
wire na142_1;
wire na143_1;
wire na144_2;
wire na145_1;
wire na146_2;
wire na147_2;
wire na148_1;
wire na149_2;
wire na150_1;
wire na151_2;
wire na152_1;
wire na153_1;
wire na154_1;
wire na155_1;
wire na155_2;
wire na158_2;
wire na159_1;
wire na160_1;
wire na160_1_i;
wire na161_1;
wire na162_1;
wire na163_1;
wire na164_1;
wire na164_1_i;
wire na165_2;
wire na166_1;
wire na166_1_i;
wire na167_1;
wire na167_1_i;
wire na167_2;
wire na167_2_i;
wire na168_1;
wire na169_1;
wire na170_1;
wire na170_1_i;
wire na171_1;
wire na171_1_i;
wire na172_1;
wire na173_2;
wire na173_2_i;
wire na175_1;
wire na176_2;
wire na177_1;
wire na177_2;
wire na178_1;
wire na179_1;
wire na179_2;
wire na180_1;
wire na181_1;
wire na182_1;
wire na182_2;
wire na184_1;
wire na184_2;
wire na186_1;
wire na187_2;
wire na188_2;
wire na189_2;
wire na190_1;
wire na191_1;
wire na192_1;
wire na193_1;
wire na193_2;
wire na194_1;
wire na195_2;
wire na196_2;
wire na198_1;
wire na199_1;
wire na200_1;
wire na201_1;
wire na202_2;
wire na203_2;
wire na204_1;
wire na206_1;
wire na207_1;
wire na208_2;
wire na209_2;
wire na210_1;
wire na211_2;
wire na212_1;
wire na213_1;
wire na214_2;
wire na215_2;
wire na216_1;
wire na217_2;
wire na218_1;
wire na218_1_i;
wire na219_1;
wire na219_1_i;
wire na219_2;
wire na219_2_i;
wire na220_2;
wire na221_1;
wire na222_1;
wire na223_2;
wire na224_1;
wire na224_1_i;
wire na225_1;
wire na226_1;
wire na227_1;
wire na227_1_i;
wire na227_2;
wire na227_2_i;
wire na228_1;
wire na229_2;
wire na229_2_i;
wire na230_1;
wire na231_1;
wire na231_1_i;
wire na231_2;
wire na231_2_i;
wire na232_1;
wire na233_1;
wire na234_1;
wire na235_1;
wire na237_1;
wire na238_1;
wire na241_1;
wire na241_1_i;
wire na242_2;
wire na244_2;
wire na244_2_i;
wire na246_1;
wire na247_1;
wire na248_2;
wire na249_1;
wire na250_2;
wire na251_1;
wire na252_2;
wire na253_1;
wire na254_2;
wire na254_2_i;
wire na255_1;
wire na256_1;
wire na256_1_i;
wire na257_1;
wire na258_1;
wire na258_1_i;
wire na259_1;
wire na260_1;
wire na260_1_i;
wire na262_1;
wire na262_2;
wire na263_1;
wire na263_1_i;
wire na263_2;
wire na263_2_i;
wire na264_1;
wire na265_1;
wire na265_1_i;
wire na266_1;
wire na267_1;
wire na267_2;
wire na269_1;
wire na270_1;
wire na270_1_i;
wire na270_2;
wire na270_2_i;
wire na271_1;
wire na272_2;
wire na272_2_i;
wire na273_2;
wire na275_1;
wire na276_1;
wire na276_1_i;
wire na281_1;
wire na282_2;
wire na282_2_i;
wire na283_1;
wire na284_1;
wire na286_2;
wire na287_1;
wire na287_1_i;
wire na288_1;
wire na288_2;
wire na289_2;
wire na290_1;
wire na291_2;
wire na291_2_i;
wire na292_1;
wire na292_1_i;
wire na293_2;
wire na293_2_i;
wire na294_2;
wire na295_1;
wire na297_1;
wire na297_1_i;
wire na297_2;
wire na297_2_i;
wire na298_1;
wire na298_1_i;
wire na299_1;
wire na299_1_i;
wire na299_2;
wire na299_2_i;
wire na300_1;
wire na300_1_i;
wire na300_2;
wire na300_2_i;
wire na304_1;
wire na306_1;
wire na308_1;
wire na309_1;
wire na309_1_i;
wire na309_2;
wire na309_2_i;
wire na311_1;
wire na311_2;
wire na312_1;
wire na314_1;
wire na314_1_i;
wire na314_2;
wire na314_2_i;
wire na315_1;
wire na316_1;
wire na316_1_i;
wire na316_2;
wire na316_2_i;
wire na317_1;
wire na318_1;
wire na318_1_i;
wire na318_2;
wire na318_2_i;
wire na319_1;
wire na321_1;
wire na322_1;
wire na322_1_i;
wire na323_1;
wire na323_1_i;
wire na323_2;
wire na323_2_i;
wire na324_2;
wire na324_2_i;
wire na325_1;
wire na328_2;
wire na328_2_i;
wire na330_2;
wire na331_1;
wire na331_1_i;
wire na332_2;
wire na333_2;
wire na334_1;
wire na335_1;
wire na335_1_i;
wire na336_1;
wire na337_1;
wire na337_1_i;
wire na337_2;
wire na337_2_i;
wire na338_2;
wire na339_1;
wire na340_2;
wire na341_1;
wire na341_1_i;
wire na342_1;
wire na343_1;
wire na343_1_i;
wire na343_2;
wire na343_2_i;
wire na344_2;
wire na345_1;
wire na346_2;
wire na347_1;
wire na347_1_i;
wire na348_1;
wire na349_1;
wire na350_2;
wire na351_1;
wire na351_1_i;
wire na352_1;
wire na353_1;
wire na353_1_i;
wire na353_2;
wire na353_2_i;
wire na354_1;
wire na355_2;
wire na355_2_i;
wire na356_2;
wire na357_1;
wire na358_2;
wire na359_2;
wire na359_2_i;
wire na360_1;
wire na362_1;
wire na363_2;
wire na364_1;
wire na365_2;
wire na365_2_i;
wire na366_1;
wire na366_2;
wire na367_1;
wire na367_1_i;
wire na367_2;
wire na367_2_i;
wire na368_1;
wire na368_1_i;
wire na369_2;
wire na370_1;
wire na371_1;
wire na371_1_i;
wire na372_1;
wire na372_1_i;
wire na374_2;
wire na375_1;
wire na375_2;
wire na376_1;
wire na377_1;
wire na377_2;
wire na378_1;
wire na379_2;
wire na379_2_i;
wire na380_1;
wire na381_1;
wire na382_1;
wire na383_1;
wire na384_1;
wire na385_2;
wire na385_2_i;
wire na386_1;
wire na388_2;
wire na388_2_i;
wire na389_2;
wire na390_1;
wire na391_1;
wire na391_1_i;
wire na391_2;
wire na391_2_i;
wire na392_1;
wire na394_1;
wire na395_1;
wire na396_1;
wire na396_1_i;
wire na397_2;
wire na397_2_i;
wire na399_2;
wire na400_2;
wire na402_1;
wire na402_1_i;
wire na402_2;
wire na402_2_i;
wire na403_1;
wire na404_1;
wire na405_1;
wire na407_2;
wire na409_2;
wire na410_1;
wire na410_1_i;
wire na411_1;
wire na412_1;
wire na412_1_i;
wire na412_2;
wire na412_2_i;
wire na413_2;
wire na415_1;
wire na416_1;
wire na416_1_i;
wire na417_2;
wire na418_2;
wire na418_2_i;
wire na419_1;
wire na420_2;
wire na420_2_i;
wire na421_1;
wire na421_1_i;
wire na421_2;
wire na421_2_i;
wire na422_1;
wire na425_1;
wire na426_1;
wire na427_1;
wire na427_1_i;
wire na427_2;
wire na427_2_i;
wire na428_1;
wire na429_1;
wire na431_1;
wire na432_1;
wire na432_1_i;
wire na432_2;
wire na432_2_i;
wire na433_1;
wire na435_1;
wire na436_1;
wire na436_1_i;
wire na436_2;
wire na436_2_i;
wire na437_1;
wire na439_1;
wire na440_1;
wire na441_2;
wire na441_2_i;
wire na442_1;
wire na443_1;
wire na446_1;
wire na448_2;
wire na449_1;
wire na450_2;
wire na451_1;
wire na451_1_i;
wire na452_1;
wire na453_2;
wire na453_2_i;
wire na454_2;
wire na456_1;
wire na456_1_i;
wire na457_2;
wire na458_2;
wire na459_2;
wire na459_2_i;
wire na460_1;
wire na461_1;
wire na461_1_i;
wire na461_2;
wire na461_2_i;
wire na462_1;
wire na464_1;
wire na465_1;
wire na465_1_i;
wire na466_1;
wire na467_1;
wire na467_1_i;
wire na468_1;
wire na468_1_i;
wire na470_1;
wire na470_2;
wire na471_1;
wire na472_2;
wire na473_2;
wire na473_2_i;
wire na474_1;
wire na475_2;
wire na476_1;
wire na477_1;
wire na477_1_i;
wire na478_1;
wire na479_1;
wire na480_1;
wire na481_1;
wire na481_1_i;
wire na482_1;
wire na483_1;
wire na484_1;
wire na485_2;
wire na485_2_i;
wire na486_1;
wire na487_2;
wire na488_1;
wire na489_2;
wire na489_2_i;
wire na490_1;
wire na491_1;
wire na492_1;
wire na493_2;
wire na494_1;
wire na494_1_i;
wire na495_1;
wire na497_2;
wire na497_2_i;
wire na498_2;
wire na498_2_i;
wire na499_1;
wire na499_1_i;
wire na499_2;
wire na499_2_i;
wire na501_1;
wire na501_1_i;
wire na501_2;
wire na501_2_i;
wire na503_1;
wire na503_1_i;
wire na503_2;
wire na503_2_i;
wire na505_1;
wire na505_1_i;
wire na505_2;
wire na505_2_i;
wire na507_1;
wire na507_1_i;
wire na507_2;
wire na507_2_i;
wire na509_1;
wire na509_1_i;
wire na509_2;
wire na509_2_i;
wire na511_1;
wire na511_1_i;
wire na511_2;
wire na511_2_i;
wire na513_1;
wire na513_1_i;
wire na513_2;
wire na513_2_i;
wire na515_1;
wire na515_1_i;
wire na515_2;
wire na515_2_i;
wire na517_1;
wire na517_1_i;
wire na517_2;
wire na517_2_i;
wire na519_1;
wire na519_1_i;
wire na519_2;
wire na519_2_i;
wire na522_1;
wire na522_1_i;
wire na523_1;
wire na523_1_i;
wire na523_2;
wire na523_2_i;
wire na525_1;
wire na525_1_i;
wire na525_2;
wire na525_2_i;
wire na526_1;
wire na527_2;
wire na528_1;
wire na529_1;
wire na529_1_i;
wire na533_1;
wire na535_1;
wire na535_2;
wire na536_1;
wire na536_2;
wire na537_1;
wire na537_1_i;
wire na541_1;
wire na543_1;
wire na543_2;
wire na544_1;
wire na544_2;
wire na545_1;
wire na546_1;
wire na547_2;
wire na548_1;
wire na549_2;
wire na550_1;
wire na551_1;
wire na552_2;
wire na553_2;
wire na554_2;
wire na555_2;
wire na556_2;
wire na557_1;
wire na558_2;
wire na559_1;
wire na560_1;
wire na576_1;
wire na577_1;
wire na578_1;
wire na578_1_i;
wire na578_2;
wire na578_2_i;
wire na579_1;
wire na580_1;
wire na581_1;
wire na581_1_i;
wire na581_2;
wire na581_2_i;
wire na582_4;
wire na583_1;
wire na583_4;
wire na604_4;
wire na608_4;
wire na610_1;
wire na614_4;
wire na615_1;
wire na615_4;
wire na636_4;
wire na640_4;
wire na642_1;
wire na648_1;
wire na648_2;
wire na648_4;
wire na650_1;
wire na650_2;
wire na650_4;
wire na652_1;
wire na652_2;
wire na652_4;
wire na654_1;
wire na654_2;
wire na654_4;
wire na656_1;
wire na656_2;
wire na656_4;
wire na657_1;
wire na657_2;
wire na657_4;
wire na659_1;
wire na659_2;
wire na659_4;
wire na661_1;
wire na661_2;
wire na661_4;
wire na663_1;
wire na663_2;
wire na666_1;
wire na666_2;
wire na666_4;
wire na668_1;
wire na668_2;
wire na668_4;
wire na670_1;
wire na670_2;
wire na670_4;
wire na672_1;
wire na672_2;
wire na672_4;
wire na673_1;
wire na673_4;
wire na675_1;
wire na675_2;
wire na675_4;
wire na677_1;
wire na677_2;
wire na677_4;
wire na679_1;
wire na679_2;
wire na679_4;
wire na681_1;
wire na681_2;
wire na681_4;
wire na683_1;
wire na683_2;
wire na684_1;
wire na684_4;
wire na685_1;
wire na685_2;
wire na685_4;
wire na687_1;
wire na687_2;
wire na687_4;
wire na689_1;
wire na690_1;
wire na690_4;
wire na691_1;
wire na691_2;
wire na691_4;
wire na693_1;
wire na693_2;
wire na693_4;
wire na695_1;
wire na695_4;
wire na696_1;
wire na697_1;
wire na697_2;
wire na697_4;
wire na699_1;
wire na699_2;
wire na699_4;
wire na701_1;
wire na702_1;
wire na702_4;
wire na703_1;
wire na703_2;
wire na703_4;
wire na705_1;
wire na705_2;
wire na705_4;
wire na707_1;
wire na707_2;
wire na709_1;
wire na709_4;
wire na711_1;
wire na711_2;
wire na711_4;
wire na713_1;
wire na713_2;
wire na713_4;
wire na715_1;
wire na715_2;
wire na715_4;
wire na717_1;
wire na717_2;
wire na717_4;
wire na719_1;
wire na719_2;
wire na719_4;
wire na720_1;
wire na720_2;
wire na720_4;
wire na722_1;
wire na722_2;
wire na722_4;
wire na724_1;
wire na724_2;
wire na724_4;
wire na726_1;
wire na726_2;
wire na726_4;
wire na728_1;
wire na730_1;
wire na730_2;
wire na730_4;
wire na732_1;
wire na732_2;
wire na732_4;
wire na734_1;
wire na734_2;
wire na734_4;
wire na736_1;
wire na736_2;
wire na736_4;
wire na737_1;
wire na737_4;
wire na739_1;
wire na739_1_i;
wire na739_2;
wire na739_4;
wire na741_1;
wire na741_1_i;
wire na741_2;
wire na741_4;
wire na743_1;
wire na743_1_i;
wire na743_2;
wire na743_4;
wire na745_1;
wire na745_1_i;
wire na745_2;
wire na745_4;
wire na747_1;
wire na747_1_i;
wire na747_2;
wire na747_4;
wire na748_1;
wire na748_1_i;
wire na748_2;
wire na748_4;
wire na750_1;
wire na750_1_i;
wire na750_2;
wire na750_4;
wire na752_1;
wire na752_1_i;
wire na752_2;
wire na755_1;
wire na755_1_i;
wire na755_2;
wire na755_4;
wire na757_1;
wire na757_1_i;
wire na757_2;
wire na757_4;
wire na759_1;
wire na759_1_i;
wire na759_2;
wire na759_4;
wire na761_1;
wire na761_1_i;
wire na761_2;
wire na761_4;
wire na762_1;
wire na762_4;
wire na764_1;
wire na764_2;
wire na764_4;
wire na766_1;
wire na766_2;
wire na766_4;
wire na768_1;
wire na768_2;
wire na768_4;
wire na770_1;
wire na770_2;
wire na770_4;
wire na772_1;
wire na772_2;
wire na773_1;
wire na773_4;
wire na774_1;
wire na774_2;
wire na774_4;
wire na776_1;
wire na776_2;
wire na776_4;
wire na778_1;
wire na779_1;
wire na779_4;
wire na780_1;
wire na780_2;
wire na780_4;
wire na782_1;
wire na782_2;
wire na782_4;
wire na784_1;
wire na784_4;
wire na785_1;
wire na786_1;
wire na786_2;
wire na786_4;
wire na788_1;
wire na788_2;
wire na788_4;
wire na790_1;
wire na790_2;
wire na790_4;
wire na792_1;
wire na793_1;
wire na793_4;
wire na794_1;
wire na794_2;
wire na794_4;
wire na796_1;
wire na796_2;
wire na796_4;
wire na798_1;
wire na798_2;
wire na798_4;
wire na800_1;
wire na801_1;
wire na801_4;
wire na803_1;
wire na803_2;
wire na803_4;
wire na805_1;
wire na805_2;
wire na805_4;
wire na807_1;
wire na807_2;
wire na807_4;
wire na809_1;
wire na809_2;
wire na809_4;
wire na811_1;
wire na811_2;
wire na811_4;
wire na812_1;
wire na812_2;
wire na812_4;
wire na814_1;
wire na814_2;
wire na814_4;
wire na816_1;
wire na816_2;
wire na816_4;
wire na818_1;
wire na818_2;
wire na818_4;
wire na820_1;
wire na822_1;
wire na822_2;
wire na822_4;
wire na824_1;
wire na824_2;
wire na824_4;
wire na826_1;
wire na826_2;
wire na826_4;
wire na828_1;
wire na828_2;
wire na828_4;
wire na829_1;
wire na829_4;
wire na831_1;
wire na831_1_i;
wire na831_2;
wire na831_4;
wire na833_1;
wire na833_1_i;
wire na833_2;
wire na833_4;
wire na835_1;
wire na835_1_i;
wire na835_2;
wire na835_4;
wire na837_1;
wire na837_1_i;
wire na837_2;
wire na837_4;
wire na839_1;
wire na839_1_i;
wire na839_2;
wire na839_4;
wire na840_1;
wire na840_1_i;
wire na840_2;
wire na840_4;
wire na842_1;
wire na842_1_i;
wire na842_2;
wire na842_4;
wire na844_1;
wire na844_1_i;
wire na844_2;
wire na847_1;
wire na847_1_i;
wire na847_2;
wire na847_4;
wire na849_1;
wire na849_1_i;
wire na849_2;
wire na849_4;
wire na851_1;
wire na851_1_i;
wire na851_2;
wire na851_4;
wire na853_1;
wire na853_1_i;
wire na853_2;
wire na853_4;
wire na900_1;
wire na900_1_i;
wire na902_2;
wire na902_2_i;
wire na906_1;
wire na906_1_i;
wire na906_2;
wire na906_2_i;
wire na908_1;
wire na908_1_i;
wire na908_2;
wire na908_2_i;
wire na912_1;
wire na912_1_i;
wire na912_2;
wire na912_2_i;
wire na916_1;
wire na916_1_i;
wire na918_2;
wire na918_2_i;
wire na920_1;
wire na920_1_i;
wire na920_2;
wire na920_2_i;
wire na922_1;
wire na922_1_i;
wire na923_2;
wire na923_2_i;
wire na924_2;
wire na924_2_i;
wire na925_2;
wire na925_2_i;
wire na926_1;
wire na926_1_i;
wire na927_2;
wire na927_2_i;
wire na928_1;
wire na928_1_i;
wire na929_2;
wire na929_2_i;
wire na993_1;
wire na993_1_i;
wire na994_1;
wire na994_1_i;
wire na994_2;
wire na994_2_i;
wire na996_1;
wire na996_1_i;
wire na996_2;
wire na996_2_i;
wire oled_dc;
wire na1010_2;
wire na1010_2_i;
wire na1012_1;
wire na1012_1_i;
wire na1016_1;
wire na1016_1_i;
wire na1016_2;
wire na1016_2_i;
wire na1018_1;
wire na1018_1_i;
wire na1018_2;
wire na1018_2_i;
wire na1022_1;
wire na1022_1_i;
wire na1022_2;
wire na1022_2_i;
wire na1026_2;
wire na1026_2_i;
wire na1028_1;
wire na1028_1_i;
wire na1030_1;
wire na1030_1_i;
wire na1030_2;
wire na1030_2_i;
wire na1032_2;
wire na1032_2_i;
wire na1033_1;
wire na1033_1_i;
wire na1034_2;
wire na1034_2_i;
wire na1035_1;
wire na1035_1_i;
wire na1036_1;
wire na1036_1_i;
wire na1037_1;
wire na1037_1_i;
wire na1038_2;
wire na1038_2_i;
wire na1039_1;
wire na1039_1_i;
wire na1115_2;
wire na1115_2_i;
wire na1116_1;
wire na1116_1_i;
wire na1116_2;
wire na1116_2_i;
wire na1118_1;
wire na1118_1_i;
wire na1118_2;
wire na1118_2_i;
wire na1122_1;
wire na1123_1;
wire na1124_1;
wire na1125_1;
wire na1126_1;
wire na1127_1;
wire na1128_1;
wire na1129_1;
wire na1130_1;
wire na1131_1;
wire na1132_1;
wire na1133_1;
wire na1133_1_i;
wire na1134_1;
wire na1135_1;
wire na1136_1;
wire na1136_1_i;
wire na1137_1;
wire na1138_1;
wire na1138_1_i;
wire na1139_1;
wire na1140_1;
wire na1141_1;
wire na1141_1_i;
wire na1142_1;
wire na1143_1;
wire na1143_1_i;
wire na1144_1;
wire na1145_1;
wire na1146_1;
wire na1146_1_i;
wire na1147_1;
wire na1147_1_i;
wire na1148_1;
wire na1149_1;
wire na1150_1;
wire na1150_1_i;
wire na1151_1;
wire na1152_1;
wire na1153_1;
wire na1154_1;
wire na1155_1;
wire na1156_1;
wire na1157_1;
wire na1158_1;
wire na1159_1;
wire na1160_1;
wire na1161_1;
wire na1162_1;
wire na1163_1;
wire na1164_1;
wire na1165_1;
wire na1166_1;
wire na1167_1;
wire na1168_1;
wire na1169_1;
wire na1170_1;
wire na1171_1;
wire na1172_1;
wire na1173_1;
wire na1174_1;
wire na1175_1;
wire na1176_1;
wire na1177_1;
wire na1178_1;
wire na1179_1;
wire na1192_3;
wire na1192_4;
wire na1192_5;
wire na1192_6;
wire na1193_1;
wire na1194_1;
wire na1194_2;
wire na1195_2;
wire na1196_1;
wire na1197_1;
wire na1197_2;
wire na1198_2;
wire na1199_1;
wire na1200_1;
wire na1201_1;
wire na1203_1;
wire na1204_2;
wire na1205_2;
wire na1206_1;
wire na1207_1;
wire na1207_4;
wire na1208_1;
wire na1208_2;
wire na1209_1;
wire na1210_1;
wire na1210_2;
wire na1212_1;
wire na1214_1;
wire na1217_1;
wire na1218_2;
wire na1219_1;
wire na1220_1;
wire na1221_1;
wire na1224_1;
wire na1225_2;
wire na1226_1;
wire na1227_2;
wire na1228_2;
wire na1229_1;
wire na1230_2;
wire na1232_1;
wire na1234_1;
wire na1236_1;
wire na1237_2;
wire na1238_1;
wire na1239_1;
wire na1240_1;
wire na1241_1;
wire na1242_1;
wire na1243_2;
wire na1244_1;
wire na1245_1;
wire na1246_1;
wire na1247_1;
wire na1248_2;
wire na1250_1;
wire na1251_2;
wire na1252_2;
wire na1253_2;
wire na1254_1;
wire na1255_2;
wire na1256_1;
wire na1257_1;
wire na1258_2;
wire na1260_2;
wire na1261_1;
wire na1264_1;
wire na1266_1;
wire na1267_1;
wire na1270_1;
wire na1271_1;
wire na1272_1;
wire na1273_2;
wire na1274_2;
wire na1275_1;
wire na1276_2;
wire na1278_1;
wire na1280_1;
wire na1281_1;
wire na1282_1;
wire na1284_1;
wire na1285_1;
wire na1286_1;
wire na1289_1;
wire na1290_1;
wire na1291_1;
wire na1292_1;
wire na1293_1;
wire na1298_1;
wire na1299_1;
wire na1300_1;
wire na1301_2;
wire na1302_1;
wire na1303_2;
wire na1304_1;
wire na1308_1;
wire na1311_2;
wire na1312_1;
wire na1313_1;
wire na1314_2;
wire na1321_1;
wire na1325_1;
wire na1327_2;
wire na1329_1;
wire na1333_1;
wire na1334_1;
wire na1335_1;
wire na1340_1;
wire na1345_1;
wire na1346_2;
wire na1347_2;
wire na1348_1;
wire na1349_2;
wire na1350_1;
wire na1351_1;
wire na1352_2;
wire na1353_1;
wire na1356_1;
wire na1357_1;
wire na1358_1;
wire na1359_1;
wire na1359_2;
wire na1360_1;
wire na1361_1;
wire na1363_1;
wire na1363_2;
wire na1364_1;
wire na1365_1;
wire na1366_1;
wire na1367_1;
wire na1370_1;
wire na1371_1;
wire na1372_1;
wire na1375_1;
wire na1378_1;
wire na1379_1;
wire na1380_2;
wire na1381_2;
wire na1382_1;
wire na1383_1;
wire na1386_1;
wire na1387_1;
wire na1388_1;
wire na1408_1;
wire na1409_2;
wire na1410_1;
wire na1411_1;
wire na1412_2;
wire na1413_2;
wire na1414_1;
wire na1415_2;
wire na1416_1;
wire na1417_1;
wire na1418_1;
wire na1419_1;
wire na1422_1;
wire na1424_1;
wire na1425_1;
wire na1426_1;
wire na1427_1;
wire na1428_1;
wire na1429_1;
wire na1430_1;
wire na1431_1;
wire na1432_1;
wire na1433_1;
wire na1434_1;
wire na1435_1;
wire na1436_1;
wire na1437_1;
wire na1438_1;
wire na1439_1;
wire na1440_1;
wire na1441_1;
wire na1441_2;
wire na1442_1;
wire na1444_1;
wire na1445_2;
wire na1447_1;
wire na1448_1;
wire na1449_1;
wire na1450_1;
wire na1451_1;
wire na1452_1;
wire na1455_1;
wire na1456_1;
wire na1457_1;
wire na1460_1;
wire na1463_1;
wire na1466_1;
wire na1469_1;
wire na1472_1;
wire na1475_1;
wire na1476_1;
wire na1478_2;
wire na1479_1;
wire na1480_1;
wire na1481_1;
wire na1482_1;
wire na1483_1;
wire na1484_2;
wire na1486_1;
wire na1487_1;
wire na1489_1;
wire na1490_1;
wire na1491_1;
wire na1492_2;
wire na1493_1;
wire na1494_1;
wire na1495_1;
wire na1496_1;
wire na1497_1;
wire na1498_1;
wire na1500_1;
wire na1501_1;
wire na1502_2;
wire na1504_1;
wire na1506_1;
wire na1507_1;
wire na1508_1;
wire na1510_1;
wire na1511_1;
wire na1514_1;
wire na1515_1;
wire na1516_1;
wire na1517_2;
wire na1518_1;
wire na1519_2;
wire na1520_1;
wire na1521_1;
wire na1522_2;
wire na1524_1;
wire na1525_2;
wire na1526_1;
wire na1527_1;
wire na1528_1;
wire na1529_1;
wire na1530_1;
wire na1531_1;
wire na1532_1;
wire na1534_2;
wire na1535_1;
wire na1537_1;
wire na1538_1;
wire na1539_2;
wire na1540_2;
wire na1541_2;
wire na1542_2;
wire na1543_2;
wire na1544_2;
wire na1545_2;
wire na1546_2;
wire na1547_2;
wire na1548_2;
wire na1549_2;
wire na1550_2;
wire na1551_2;
wire na1552_2;
wire na1553_2;
wire na1554_2;
wire na1555_2;
wire na1556_2;
wire na1557_2;
wire na1558_2;
wire na1559_2;
wire na1560_2;
wire na1561_2;
wire na1562_2;
wire na1563_2;
wire na1564_2;
wire na1565_2;
wire na1566_2;
wire na1567_2;
wire na1568_2;
wire na1569_2;
wire na1570_2;
wire na1571_2;
wire na1572_2;
wire na1573_2;
wire na1574_2;
wire na1575_2;
wire na1576_2;
wire na1577_2;
wire na1578_2;
wire na1579_2;
wire na1580_2;
wire na1581_2;
wire na1582_2;
wire na1583_2;
wire na1584_2;
wire na1585_2;
wire na1586_2;
wire na1587_2;
wire na1588_2;
wire na1589_2;
wire na1590_2;
wire na1591_2;
wire na1592_2;
wire na1593_2;
wire na1594_2;
wire na1595_2;
wire na1596_2;
wire na1597_2;
wire na1598_2;
wire na1599_2;
wire na1600_2;
wire na1601_2;
wire na1602_2;
wire na1603_2;
wire na1604_2;
wire na1605_2;
wire na1606_2;
wire na1607_2;
wire na1608_2;
wire na1609_2;
wire na1610_2;
wire na1611_2;
wire na1612_2;
wire na1613_2;
wire na1614_2;
wire na1615_2;
wire na1616_2;
wire na1617_2;
wire na1618_2;
wire na1619_2;
wire na1620_2;
wire na1621_2;
wire na1622_2;
wire na1623_2;
wire na1624_2;
wire na1625_2;
wire na1626_2;
wire na1627_2;
wire na1628_2;
wire na1629_2;
wire na1630_2;
wire na1631_2;
wire na1632_2;
wire na1633_2;
wire na1634_2;
wire na1635_2;
wire na1636_2;
wire na1637_2;
wire na1638_2;
wire na1639_2;
wire na1640_2;
wire na1641_2;
wire na1642_2;
wire na1643_2;
wire na1644_2;
wire na1645_2;
wire na1646_2;
wire na1647_2;
wire na1648_2;
wire na1649_2;
wire na1650_2;
wire na1651_2;
wire na1652_2;
wire na1653_2;
wire na1654_2;
wire na1655_2;
wire na1656_2;
wire na1657_2;
wire na1658_2;
wire na1659_2;
wire na1660_2;
wire na1661_2;
wire na1662_2;
wire na1663_2;
wire na1664_2;
wire na1665_2;
wire na1666_2;
wire na1667_2;
wire na1668_2;
wire na1669_2;
wire na1670_2;
wire na1671_2;
wire na1672_2;
wire na1673_2;
wire na1674_2;
wire na1675_2;
wire na1676_2;
wire na1677_2;
wire na1678_2;
wire na1679_2;
wire na1680_2;
wire na1681_2;
wire na1682_2;
wire na1683_2;
wire na1684_2;
wire na1685_2;
wire na1686_2;
wire na1687_2;
wire na1688_2;
wire na1689_2;
wire na1690_2;
wire na1691_2;
wire na1692_2;
wire na1693_2;
wire na1694_2;
wire na1695_2;
wire na1696_2;
wire na1697_2;
wire na1698_2;
wire na1699_2;
wire na1700_2;
wire na1701_2;
wire na1702_2;
wire na1703_2;
wire na1704_2;
wire na1705_2;
wire na1706_2;
wire na1707_2;
wire na1708_2;
wire oled_clk;
wire oled_csn;
wire na1539_10;
wire na1540_10;
wire na1541_10;
wire na1542_10;
wire na1543_10;
wire na1544_10;
wire na1545_10;
wire na1546_10;
wire na1547_10;
wire na1548_10;
wire oled_dc_1;
wire oled_mosi;
wire oled_resn;
wire oled_clk_1;
wire oled_mosi_1;
wire oled_resn_1;

// C_///OR/      x32y106     80'h00_0060_00_0000_0C0E_FF0D
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1_4 ( .OUT(na1_2), .IN1(~na610_1), .IN2(na1193_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x42y104     80'h00_0018_00_0000_0888_FDAB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a6_1 ( .OUT(na6_1), .IN1(na780_1), .IN2(~na219_1), .IN3(na1200_1), .IN4(1'b0), .IN5(~na785_1), .IN6(na219_2), .IN7(1'b1),
                   .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x40y104     80'h00_0018_00_0000_0C88_DBFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a7_1 ( .OUT(na7_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na780_1), .IN6(~na219_1), .IN7(~na1682_2), .IN8(na1608_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x33y105     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a8_4 ( .OUT(na8_2), .IN1(~na10_1), .IN2(1'b0), .IN3(~na276_1), .IN4(na1_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y105     80'h00_0018_00_0000_0888_8841
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a10_1 ( .OUT(na10_1), .IN1(~na1199_1), .IN2(~na1618_2), .IN3(~na1196_1), .IN4(na6_1), .IN5(na1195_2), .IN6(na1194_1), .IN7(na1702_2),
                    .IN8(na1198_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x42y108     80'h00_FE18_00_0000_0888_FC3F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a11_1 ( .OUT(na11_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na12_1), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a11_5 ( .OUT(na11_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na11_1) );
// C_MX2b////      x36y106     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na13_1), .IN5(~na683_1), .IN6(1'b0), .IN7(~na1549_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x44y104     80'h00_0078_00_0000_0C88_5AC3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na265_1), .IN6(1'b1), .IN7(~na14_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a13_4 ( .OUT(na13_2), .IN1(1'b1), .IN2(~na32_1), .IN3(1'b1), .IN4(na420_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x40y111     80'h00_0018_00_0000_0888_281C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a14_1 ( .OUT(na14_1), .IN1(1'b1), .IN2(na184_2), .IN3(~na179_2), .IN4(~na11_2), .IN5(na182_2), .IN6(na1554_2), .IN7(na17_2),
                    .IN8(~na177_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////D      x32y115     80'h00_FE18_00_0000_0888_FFDC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a17_1 ( .OUT(na17_1), .IN1(1'b0), .IN2(na470_2), .IN3(~na1203_1), .IN4(na1204_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a17_5 ( .OUT(na17_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na17_1) );
// C_ORAND////D      x42y112     80'h00_FE18_00_0000_0888_FFDC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a19_1 ( .OUT(na19_1), .IN1(1'b0), .IN2(na470_2), .IN3(~na1205_2), .IN4(na1206_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a19_5 ( .OUT(na19_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na19_1) );
// C_///ORAND/      x45y118     80'h00_0060_00_0000_0C08_FF7B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a20_4 ( .OUT(na20_2), .IN1(na265_1), .IN2(~na1554_2), .IN3(~na1658_2), .IN4(~na13_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x41y113     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a21_1 ( .OUT(na21_1), .IN1(1'b1), .IN2(na20_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na17_1), .IN8(na11_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x29y103     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1), .IN1(1'b1), .IN2(~na1621_2), .IN3(1'b0), .IN4(1'b0), .IN5(na23_1), .IN6(na371_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y109     80'h00_0018_00_0000_0888_3313
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a23_1 ( .OUT(na23_1), .IN1(1'b1), .IN2(~na219_1), .IN3(~na272_2), .IN4(~na270_2), .IN5(1'b1), .IN6(~na219_2), .IN7(1'b1),
                    .IN8(~na270_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x42y101     80'h00_0018_00_0000_0CEE_C300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a25_1 ( .OUT(na25_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na642_1), .IN7(1'b0), .IN8(na30_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x41y106     80'h00_0018_00_0040_0AC4_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a29_1 ( .OUT(na29_1), .IN1(~na397_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na25_1), .IN8(na30_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x40y108     80'h00_0018_00_0000_0888_A8A8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a30_1 ( .OUT(na30_1), .IN1(na1209_1), .IN2(na1210_1), .IN3(na1208_2), .IN4(1'b1), .IN5(na1212_1), .IN6(na1210_2), .IN7(na1208_1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x43y89     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a31_1 ( .OUT(na31_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na420_2), .IN5(1'b0), .IN6(na32_1), .IN7(1'b0), .IN8(na1649_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x41y92     80'h00_0018_00_0000_0888_31F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a32_1 ( .OUT(na32_1), .IN1(~na402_2), .IN2(~na1643_2), .IN3(1'b1), .IN4(1'b1), .IN5(~na402_1), .IN6(~na410_1), .IN7(1'b1),
                    .IN8(~na1644_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x37y109     80'h00_0018_00_0000_0C88_7BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a35_1 ( .OUT(na35_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na23_1), .IN6(~na1122_1), .IN7(~na1681_2), .IN8(~na36_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x36y112     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1217_1), .IN6(na1556_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y103     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a39_4 ( .OUT(na39_2), .IN1(na1363_2), .IN2(1'b1), .IN3(1'b1), .IN4(na292_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x32y99     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a44_1 ( .OUT(na44_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1178_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na537_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x43y88     80'h00_0078_00_0000_0C88_5A28
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a48_1 ( .OUT(na48_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na707_2), .IN6(1'b1), .IN7(~na49_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a48_4 ( .OUT(na48_2), .IN1(na467_1), .IN2(na1441_2), .IN3(na1551_2), .IN4(~na420_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x44y85     80'h00_0018_00_0000_0888_A884
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a49_1 ( .OUT(na49_1), .IN1(~na135_1), .IN2(na1634_2), .IN3(na497_2), .IN4(na343_2), .IN5(na135_2), .IN6(na337_2), .IN7(na1633_2),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x33y96     80'h00_FE00_80_0000_0C88_ACAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a51_1 ( .OUT(na51_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1221_1), .IN7(na44_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a51_2 ( .OUT(na51_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na51_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a51_4 ( .OUT(na51_2_i), .IN1(na1286_1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a51_5 ( .OUT(na51_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na51_2_i) );
// C_MX2b////      x32y102     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a54_1 ( .OUT(na54_1), .IN1(1'b1), .IN2(1'b1), .IN3(na55_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na256_1), .IN7(1'b0), .IN8(~na1_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x30y105     80'h00_0018_00_0000_0C88_4AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1363_2), .IN6(1'b1), .IN7(~na1555_2), .IN8(na292_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x25y93     80'h00_0018_00_0000_0888_4841
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a56_1 ( .OUT(na56_1), .IN1(~na258_1), .IN2(~na377_2), .IN3(~na141_2), .IN4(na1615_2), .IN5(na137_2), .IN6(na1569_2), .IN7(~na375_2),
                    .IN8(na155_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x23y88     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a57_4 ( .OUT(na57_2), .IN1(1'b1), .IN2(na256_1), .IN3(~na1219_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x33y93     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a58_1 ( .OUT(na58_1), .IN1(1'b1), .IN2(~na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1224_1), .IN8(~na811_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y94     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a61_1 ( .OUT(na61_1), .IN1(1'b1), .IN2(na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na814_1), .IN8(~na1227_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x30y92     80'h00_0018_00_0040_0A50_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a62_1 ( .OUT(na62_1), .IN1(na166_1), .IN2(1'b1), .IN3(~na1580_2), .IN4(1'b1), .IN5(na1228_2), .IN6(1'b0), .IN7(na167_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x40y97     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a63_1 ( .OUT(na63_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1229_1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a63_2 ( .OUT(na63_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na63_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a63_4 ( .OUT(na63_2_i), .IN1(na1558_2), .IN2(1'b1), .IN3(na1226_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a63_5 ( .OUT(na63_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na63_2_i) );
// C_MX2b////      x35y95     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a64_1 ( .OUT(na64_1), .IN1(1'b1), .IN2(na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na814_2), .IN8(~na1230_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x50y98     80'h00_FE00_00_0000_0CEE_C300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a66_1 ( .OUT(na66_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na470_2), .IN7(1'b0), .IN8(na1232_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a66_2 ( .OUT(na66_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na66_1_i) );
// C_///AND/      x43y99     80'h00_0060_00_0000_0C08_FF41
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a69_4 ( .OUT(na69_2), .IN1(~na397_2), .IN2(~na32_1), .IN3(~na25_1), .IN4(na420_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x44y100     80'h00_0018_00_0000_0888_BFCC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a70_1 ( .OUT(na70_1), .IN1(1'b0), .IN2(na1441_2), .IN3(1'b0), .IN4(na13_1), .IN5(1'b1), .IN6(1'b1), .IN7(na25_1), .IN8(~na13_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y107     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a72_1 ( .OUT(na72_1), .IN1(~na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1236_1), .IN8(~na734_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y118     80'h00_0018_00_0040_0A50_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a73_1 ( .OUT(na73_1), .IN1(na1141_1), .IN2(1'b1), .IN3(na1697_2), .IN4(1'b1), .IN5(na1237_2), .IN6(1'b0), .IN7(na1133_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/D      x40y85     80'h00_FE00_80_0000_0C0E_FFD0
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a74_4 ( .OUT(na74_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na44_1), .IN4(na1238_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a74_5 ( .OUT(na74_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na74_2_i) );
// C_MX2b////      x35y87     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1), .IN1(1'b1), .IN2(~na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1239_1), .IN8(~na822_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x31y87     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a77_1 ( .OUT(na77_1), .IN1(1'b1), .IN2(na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na824_1), .IN8(~na1241_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x33y88     80'h00_FE00_80_0000_0C88_ACAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1242_1), .IN7(na44_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_2 ( .OUT(na78_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a78_4 ( .OUT(na78_2_i), .IN1(na1240_1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a78_5 ( .OUT(na78_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_2_i) );
// C_MX2b////      x31y85     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a79_1 ( .OUT(na79_1), .IN1(1'b1), .IN2(na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na824_2), .IN8(~na1243_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x50y97     80'h00_FE00_80_0000_0C88_F8CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1244_1), .IN6(na470_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_2 ( .OUT(na80_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na80_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a80_4 ( .OUT(na80_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(1'b1), .IN4(na1272_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a80_5 ( .OUT(na80_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na80_2_i) );
// C_MX2b////      x50y108     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a81_1 ( .OUT(na81_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na732_2), .IN8(~na1245_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x44y90     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a83_4 ( .OUT(na83_2_i), .IN1(na1247_1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a83_5 ( .OUT(na83_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na83_2_i) );
// C_MX2b////      x34y87     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a84_1 ( .OUT(na84_1), .IN1(1'b1), .IN2(~na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1248_2), .IN8(~na826_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x28y92     80'h00_0018_00_0040_0AAF_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a85_1 ( .OUT(na85_1), .IN1(1'b1), .IN2(~na160_1), .IN3(~na1583_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na1703_2), .IN7(1'b1),
                    .IN8(~na164_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y90     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a87_1 ( .OUT(na87_1), .IN1(1'b1), .IN2(na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na828_1), .IN8(~na1251_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x29y92     80'h00_0018_00_0040_0CD6_3500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a88_1 ( .OUT(na88_1), .IN1(1'b1), .IN2(na1253_2), .IN3(~na1252_2), .IN4(1'b1), .IN5(~na166_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na164_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x38y90     80'h00_FE00_80_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1254_1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_2 ( .OUT(na89_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a89_4 ( .OUT(na89_2_i), .IN1(1'b1), .IN2(na1250_1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a89_5 ( .OUT(na89_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_2_i) );
// C_MX2b////      x35y90     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1615_2), .IN5(~na1255_2), .IN6(1'b0), .IN7(~na828_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x39y93     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a92_4 ( .OUT(na92_2_i), .IN1(na1558_2), .IN2(1'b1), .IN3(na1257_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a92_5 ( .OUT(na92_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na92_2_i) );
// C_MX2b////      x37y94     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_1 ( .OUT(na93_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1615_2), .IN5(1'b0), .IN6(~na1258_2), .IN7(1'b0), .IN8(~na803_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x27y96     80'h00_0018_00_0040_0A60_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a94_1 ( .OUT(na94_1), .IN1(na166_1), .IN2(1'b1), .IN3(1'b1), .IN4(na164_1), .IN5(1'b0), .IN6(na1253_2), .IN7(na1260_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x39y92     80'h00_FE00_00_0000_0CEE_5C00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a95_1 ( .OUT(na95_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1261_1), .IN7(~na44_1), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a95_2 ( .OUT(na95_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na95_1_i) );
// C_ORAND///ORAND/      x40y92     80'h00_0078_00_0000_0C88_5DCB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a96_1 ( .OUT(na96_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1686_2), .IN6(na256_1), .IN7(~na97_1), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a96_4 ( .OUT(na96_2), .IN1(na1617_2), .IN2(~na57_2), .IN3(1'b0), .IN4(na54_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x34y91     80'h00_0018_00_0000_0C88_23FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a97_1 ( .OUT(na97_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1225_2), .IN7(na98_2), .IN8(~na1579_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x34y91     80'h00_0060_00_0000_0C08_FF58
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a98_4 ( .OUT(na98_2), .IN1(na166_1), .IN2(na256_1), .IN3(~na167_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x37y89     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a99_4 ( .OUT(na99_2_i), .IN1(1'b1), .IN2(na1264_1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a99_5 ( .OUT(na99_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na99_2_i) );
// C_ORAND////      x35y92     80'h00_0018_00_0000_0C88_7DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a100_1 ( .OUT(na100_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1687_2), .IN6(na256_1), .IN7(~na98_2), .IN8(~na1266_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x38y94     80'h00_FE00_00_0000_0CEE_5A00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a102_1 ( .OUT(na102_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1267_1), .IN6(1'b0), .IN7(~na44_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a102_2 ( .OUT(na102_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na102_1_i) );
// C_ORAND////      x32y87     80'h00_0018_00_0000_0C88_5DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_1 ( .OUT(na103_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1688_2), .IN6(na256_1), .IN7(~na104_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x32y89     80'h00_0018_00_0000_0C88_83FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a104_1 ( .OUT(na104_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1225_2), .IN7(na98_2), .IN8(na1579_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x34y85     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a106_1 ( .OUT(na106_1), .IN1(1'b1), .IN2(na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na812_1), .IN8(~na1271_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y97     80'h00_0060_00_0000_0C08_FF21
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a107_4 ( .OUT(na107_2), .IN1(~na166_1), .IN2(~na160_1), .IN3(na167_2), .IN4(~na164_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y106     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a109_1 ( .OUT(na109_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na732_1), .IN8(~na1273_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x47y116     80'h00_0018_00_0040_0C05_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a110_1 ( .OUT(na110_1), .IN1(na1704_2), .IN2(1'b0), .IN3(na1133_1), .IN4(1'b0), .IN5(na1141_1), .IN6(1'b1), .IN7(~na1697_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/D      x50y98     80'h00_FE00_80_0000_0C0E_FF5C
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a111_4 ( .OUT(na111_2_i), .IN1(1'b0), .IN2(na1275_1), .IN3(~na1650_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a111_5 ( .OUT(na111_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na111_2_i) );
// C_MX2b////      x46y107     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a112_1 ( .OUT(na112_1), .IN1(~na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1276_2), .IN8(~na730_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x35y91     80'h00_0018_00_0000_0C88_7DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a115_1 ( .OUT(na115_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1689_2), .IN6(na256_1), .IN7(~na98_2), .IN8(~na1280_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x35y96     80'h00_FE00_00_0000_0CEE_D000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a117_1 ( .OUT(na117_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na44_1), .IN8(na1281_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a117_2 ( .OUT(na117_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na117_1_i) );
// C_MX2b////      x33y95     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a118_1 ( .OUT(na118_1), .IN1(1'b1), .IN2(na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na809_1), .IN8(na119_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x32y96     80'h00_0018_00_0040_0A55_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a119_1 ( .OUT(na119_1), .IN1(1'b0), .IN2(1'b0), .IN3(na167_1), .IN4(1'b1), .IN5(~na1282_1), .IN6(1'b0), .IN7(~na107_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x40y98     80'h00_FE00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a121_4 ( .OUT(na121_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na44_1), .IN4(na1284_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a121_5 ( .OUT(na121_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na121_2_i) );
// C_MX2b////      x34y93     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a122_1 ( .OUT(na122_1), .IN1(1'b1), .IN2(na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na809_2), .IN8(na123_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x28y96     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a123_1 ( .OUT(na123_1), .IN1(1'b1), .IN2(~na1584_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na125_2), .IN6(~na1285_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x23y93     80'h00_0060_00_0000_0C08_FF14
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a125_4 ( .OUT(na125_2), .IN1(~na166_1), .IN2(na160_1), .IN3(~na167_2), .IN4(~na164_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x31y95     80'h00_0018_00_0000_0888_FD55
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a127_1 ( .OUT(na127_1), .IN1(~na128_1), .IN2(1'b0), .IN3(~na130_1), .IN4(1'b0), .IN5(~na1690_2), .IN6(na256_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y95     80'h00_0018_00_0000_0888_F42C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1), .IN1(1'b1), .IN2(na1253_2), .IN3(na167_1), .IN4(~na164_1), .IN5(~na166_1), .IN6(na256_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x30y95     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a130_1 ( .OUT(na130_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1585_2), .IN6(na160_1), .IN7(na98_2), .IN8(na164_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x40y86     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a131_1 ( .OUT(na131_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1558_2), .IN6(1'b1), .IN7(na1289_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a131_2 ( .OUT(na131_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na131_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a131_4 ( .OUT(na131_2_i), .IN1(na1270_1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a131_5 ( .OUT(na131_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na131_2_i) );
// C_MX2b////      x36y85     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a132_1 ( .OUT(na132_1), .IN1(1'b1), .IN2(na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na812_2), .IN8(~na1290_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x39y86     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a133_1 ( .OUT(na133_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na44_1), .IN8(na1291_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a133_2 ( .OUT(na133_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na133_1_i) );
// C_MX2b////      x33y85     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a134_1 ( .OUT(na134_1), .IN1(1'b1), .IN2(~na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1292_1), .IN8(~na822_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x41y89     80'h00_FE00_80_0000_0C88_CCF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a135_1 ( .OUT(na135_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1), .IN8(na1293_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a135_2 ( .OUT(na135_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na135_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a135_4 ( .OUT(na135_2_i), .IN1(na1220_1), .IN2(na470_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a135_5 ( .OUT(na135_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na135_2_i) );
// C_///AND/      x45y94     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a136_4 ( .OUT(na136_2), .IN1(na707_1), .IN2(1'b1), .IN3(~na49_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x25y87     80'h00_FE18_00_0000_0888_3FAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a137_1 ( .OUT(na137_1), .IN1(1'b1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na138_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a137_5 ( .OUT(na137_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na137_1) );
// C_ORAND///ORAND/      x30y88     80'h00_0078_00_0000_0C88_7D7D
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na137_2), .IN6(na256_1), .IN7(~na768_1), .IN8(~na1561_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a138_4 ( .OUT(na138_2), .IN1(~na1568_2), .IN2(na256_1), .IN3(~na1560_2), .IN4(~na766_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x24y88     80'h00_FE18_00_0000_0888_3FAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a139_1 ( .OUT(na139_1), .IN1(1'b1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na138_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a139_5 ( .OUT(na139_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na139_1) );
// C_AND////D      x30y87     80'h00_FE18_00_0000_0888_AF5F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a141_1 ( .OUT(na141_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na142_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a141_5 ( .OUT(na141_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na141_1) );
// C_MX2b////      x28y85     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a142_1 ( .OUT(na142_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na768_2), .IN8(~na1570_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x25y90     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a143_1 ( .OUT(na143_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1558_2), .IN6(1'b1), .IN7(na1298_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x19y88     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a144_4 ( .OUT(na144_2), .IN1(1'b1), .IN2(na1565_2), .IN3(1'b1), .IN4(na139_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x26y87     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a145_1 ( .OUT(na145_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na137_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na139_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x24y87     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a146_4 ( .OUT(na146_2), .IN1(1'b1), .IN2(na144_2), .IN3(na142_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x26y89     80'h00_0060_00_0000_0C08_FF83
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a147_4 ( .OUT(na147_2), .IN1(1'b1), .IN2(~na1565_2), .IN3(na142_1), .IN4(na139_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x22y88     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a148_1 ( .OUT(na148_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na144_2), .IN7(~na142_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x22y88     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a149_4 ( .OUT(na149_2), .IN1(1'b1), .IN2(na150_1), .IN3(1'b1), .IN4(~na138_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x23y88     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a150_1 ( .OUT(na150_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na141_1), .IN8(~na138_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y88     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a151_4 ( .OUT(na151_2), .IN1(1'b1), .IN2(1'b1), .IN3(na44_1), .IN4(na1299_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y89     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a152_1 ( .OUT(na152_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1300_1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x27y88     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a153_1 ( .OUT(na153_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na137_1), .IN6(1'b1), .IN7(na142_1), .IN8(na138_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x28y89     80'h00_0018_00_0040_0C8C_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a154_1 ( .OUT(na154_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1705_2), .IN4(~na138_1), .IN5(1'b1), .IN6(na1566_2), .IN7(na44_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////D      x26y96     80'h00_FE18_00_0000_0888_FFAB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a155_1 ( .OUT(na155_1), .IN1(na1303_2), .IN2(~na1302_1), .IN3(na44_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a155_5 ( .OUT(na155_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na155_1) );
// C_///AND/      x26y85     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a158_4 ( .OUT(na158_2), .IN1(~na137_1), .IN2(~na150_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x23y85     80'h00_0018_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a159_1 ( .OUT(na159_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na142_1), .IN4(1'b1), .IN5(na137_1), .IN6(1'b0), .IN7(na1574_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x27y92     80'h00_FE00_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a160_1 ( .OUT(na160_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na155_1), .IN5(1'b0), .IN6(na1304_1), .IN7(1'b0), .IN8(na1124_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a160_2 ( .OUT(na160_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na160_1_i) );
// C_ORAND////      x29y87     80'h00_0018_00_0000_0C88_75FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a161_1 ( .OUT(na161_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na137_1), .IN6(1'b0), .IN7(~na141_1), .IN8(~na138_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x26y88     80'h00_0018_00_0000_0C88_BCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a162_1 ( .OUT(na162_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na1567_2), .IN7(na142_1), .IN8(~na138_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x26y85     80'h00_0018_00_0000_0CEE_CC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a163_1 ( .OUT(na163_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na153_1), .IN7(1'b0), .IN8(na148_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x26y94     80'h00_FE00_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a164_1 ( .OUT(na164_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na155_1), .IN5(1'b0), .IN6(na1125_1), .IN7(1'b0), .IN8(na138_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a164_2 ( .OUT(na164_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na164_1_i) );
// C_///AND/      x19y89     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a165_4 ( .OUT(na165_2), .IN1(1'b1), .IN2(1'b1), .IN3(na44_1), .IN4(na1308_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x27y93     80'h00_FE00_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a166_1 ( .OUT(na166_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na155_1), .IN5(1'b0), .IN6(na1126_1), .IN7(1'b0), .IN8(na138_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a166_2 ( .OUT(na166_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na166_1_i) );
// C_AND/D//AND/D      x28y95     80'h00_FE00_80_0000_0C88_3C2F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a167_1 ( .OUT(na167_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1127_1), .IN7(1'b1), .IN8(~na155_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a167_2 ( .OUT(na167_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na167_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a167_4 ( .OUT(na167_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1123_1), .IN4(~na155_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a167_5 ( .OUT(na167_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na167_2_i) );
// C_ICOMP////      x28y87     80'h00_0018_00_0000_0888_6FAC
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a168_1 ( .OUT(na168_1), .IN1(1'b0), .IN2(~na1565_2), .IN3(~na44_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na142_1), .IN8(~na138_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x27y91     80'h00_0018_00_0040_0CC1_5300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a169_1 ( .OUT(na169_1), .IN1(na1301_2), .IN2(1'b0), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1566_2), .IN7(~na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x25y97     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a170_1 ( .OUT(na170_1_i), .IN1(1'b1), .IN2(na1578_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1128_1), .IN6(na1311_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a170_2 ( .OUT(na170_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na170_1_i) );
// C_AND/D///      x27y98     80'h00_FE00_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a171_1 ( .OUT(na171_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1129_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na155_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a171_2 ( .OUT(na171_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na171_1_i) );
// C_AND////      x27y89     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a172_1 ( .OUT(na172_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1312_1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x27y98     80'h00_FE00_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a173_4 ( .OUT(na173_2_i), .IN1(1'b1), .IN2(na1130_1), .IN3(1'b1), .IN4(~na155_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a173_5 ( .OUT(na173_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na173_2_i) );
// C_MX2b////      x31y97     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a175_1 ( .OUT(na175_1), .IN1(1'b1), .IN2(na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na818_1), .IN8(~na1314_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x30y113     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a176_4 ( .OUT(na176_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na179_1), .IN4(~na177_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x30y114     80'h00_FE18_00_0000_0888_FC3F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a177_1 ( .OUT(na177_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na178_1), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a177_5 ( .OUT(na177_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na177_1) );
// C_MX2b////      x34y116     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a178_1 ( .OUT(na178_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na13_1), .IN5(1'b0), .IN6(~na677_2), .IN7(1'b0), .IN8(~na177_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x38y111     80'h00_FE18_00_0000_0888_FC5F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a179_1 ( .OUT(na179_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na180_1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a179_5 ( .OUT(na179_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na179_1) );
// C_MX2b////      x32y113     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a180_1 ( .OUT(na180_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na13_1), .IN5(~na679_2), .IN6(1'b0), .IN7(~na179_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x27y118     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a181_1 ( .OUT(na181_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na182_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na177_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x33y113     80'h00_FE18_00_0000_0888_FFF4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_1 ( .OUT(na182_1), .IN1(~na189_2), .IN2(na470_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a182_5 ( .OUT(na182_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na182_1) );
// C_AND////D      x31y116     80'h00_FE18_00_0000_0888_F3FC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a184_1 ( .OUT(na184_1), .IN1(1'b1), .IN2(na470_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na206_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a184_5 ( .OUT(na184_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na184_1) );
// C_ORAND////      x37y115     80'h00_0018_00_0000_0C88_37FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a186_1 ( .OUT(na186_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na189_2), .IN6(~na1594_2), .IN7(1'b0), .IN8(~na1593_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x37y110     80'h00_0060_00_0000_0C08_FF3B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a187_4 ( .OUT(na187_2), .IN1(na1321_1), .IN2(~na470_2), .IN3(1'b0), .IN4(~na1592_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x38y117     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a188_4 ( .OUT(na188_2), .IN1(1'b1), .IN2(na184_1), .IN3(1'b1), .IN4(na178_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x35y113     80'h00_0060_00_0000_0C08_FF7B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a189_4 ( .OUT(na189_2), .IN1(na265_1), .IN2(~na1591_2), .IN3(~na1655_2), .IN4(~na13_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x40y114     80'h00_0018_00_0000_0888_6FAC
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a190_1 ( .OUT(na190_1), .IN1(1'b0), .IN2(~na470_2), .IN3(~na1595_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na180_1), .IN8(~na178_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x42y115     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a191_1 ( .OUT(na191_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1588_2), .IN6(~na184_1), .IN7(1'b0), .IN8(~na177_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y117     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a192_1 ( .OUT(na192_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na182_1), .IN6(1'b1), .IN7(1'b1), .IN8(na178_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x30y118     80'h00_0078_00_0000_0C88_8A4C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a193_1 ( .OUT(na193_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na182_1), .IN6(1'b1), .IN7(na180_1), .IN8(na178_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a193_4 ( .OUT(na193_2), .IN1(1'b1), .IN2(na470_2), .IN3(~na180_1), .IN4(na178_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x38y118     80'h00_0018_00_0040_0AA2_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a194_1 ( .OUT(na194_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na17_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1325_1), .IN7(1'b0), .IN8(na193_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x36y114     80'h00_0060_00_0000_0C08_FFC4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a195_4 ( .OUT(na195_2), .IN1(~na189_2), .IN2(na184_1), .IN3(1'b1), .IN4(na178_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x30y116     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a196_4 ( .OUT(na196_2), .IN1(1'b1), .IN2(~na1599_2), .IN3(1'b1), .IN4(~na193_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x36y115     80'h00_0018_00_0000_0C88_BCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a198_1 ( .OUT(na198_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na470_2), .IN7(na1327_2), .IN8(~na178_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y117     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a199_1 ( .OUT(na199_1), .IN1(1'b1), .IN2(~na184_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na198_1), .IN8(~na196_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x33y116     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a200_1 ( .OUT(na200_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1597_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na190_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y114     80'h00_0018_00_0000_0C88_44FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a201_1 ( .OUT(na201_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na189_2), .IN6(na470_2), .IN7(~na180_1), .IN8(na178_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y117     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a202_4 ( .OUT(na202_2), .IN1(na189_2), .IN2(1'b1), .IN3(1'b1), .IN4(na193_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x39y113     80'h00_0060_00_0000_0C08_FF82
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a203_4 ( .OUT(na203_2), .IN1(na182_1), .IN2(~na184_1), .IN3(na180_1), .IN4(na178_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x39y116     80'h00_0018_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a204_1 ( .OUT(na204_1), .IN1(1'b0), .IN2(1'b0), .IN3(na17_1), .IN4(1'b1), .IN5(na203_2), .IN6(1'b0), .IN7(na1329_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x41y112     80'h00_0018_00_0000_0C88_7BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a206_1 ( .OUT(na206_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na265_1), .IN6(~na184_2), .IN7(~na1656_2), .IN8(~na13_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x40y116     80'h00_0018_00_0040_0C29_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a207_1 ( .OUT(na207_1), .IN1(na189_2), .IN2(1'b1), .IN3(1'b0), .IN4(na193_1), .IN5(1'b1), .IN6(~na184_1), .IN7(1'b1), .IN8(~na193_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x40y115     80'h00_0060_00_0000_0C08_FFBC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a208_4 ( .OUT(na208_2), .IN1(1'b0), .IN2(na470_2), .IN3(na1333_1), .IN4(~na178_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x42y115     80'h00_0060_00_0000_0C08_FF53
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a209_4 ( .OUT(na209_2), .IN1(1'b1), .IN2(~na184_1), .IN3(~na208_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x32y114     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a210_1 ( .OUT(na210_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na192_1), .IN6(1'b1), .IN7(~na188_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x37y113     80'h00_0060_00_0000_0C0E_FF5C
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a211_4 ( .OUT(na211_2), .IN1(1'b0), .IN2(na1334_1), .IN3(~na1650_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x44y109     80'h00_0018_00_0000_0888_7CAB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a212_1 ( .OUT(na212_1), .IN1(na265_1), .IN2(~na1553_2), .IN3(na1604_2), .IN4(1'b0), .IN5(1'b0), .IN6(na184_1), .IN7(~na1657_2),
                     .IN8(~na13_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x38y116     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a213_1 ( .OUT(na213_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1335_1), .IN6(1'b1), .IN7(na1596_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x40y110     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a214_4 ( .OUT(na214_2), .IN1(na211_2), .IN2(~na184_1), .IN3(~na198_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x32y114     80'h00_0060_00_0000_0C0E_FFCA
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a215_4 ( .OUT(na215_2), .IN1(na202_2), .IN2(1'b0), .IN3(1'b0), .IN4(na193_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x38y115     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a216_1 ( .OUT(na216_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na211_2), .IN6(~na201_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x33y115     80'h00_0060_00_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a217_4 ( .OUT(na217_2), .IN1(~na211_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na193_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x21y85     80'h00_FE00_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a218_1 ( .OUT(na218_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na218_1), .IN6(na57_2), .IN7(na44_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a218_2 ( .OUT(na218_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na218_1_i) );
// C_AND/D//AND/D      x35y106     80'h00_FE00_80_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a219_1 ( .OUT(na219_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1340_1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a219_2 ( .OUT(na219_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na219_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a219_4 ( .OUT(na219_2_i), .IN1(1'b1), .IN2(na1214_1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a219_5 ( .OUT(na219_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na219_2_i) );
// C_///ORAND/      x39y107     80'h00_0060_00_0000_0C08_FF7B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a220_4 ( .OUT(na220_2), .IN1(na23_1), .IN2(~na1151_1), .IN3(~na1675_2), .IN4(~na36_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x39y118     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a221_1 ( .OUT(na221_1), .IN1(1'b1), .IN2(na184_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na208_2), .IN8(na178_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y118     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a222_1 ( .OUT(na222_1), .IN1(1'b1), .IN2(na184_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na216_1), .IN8(na178_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x38y115     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a223_4 ( .OUT(na223_2), .IN1(1'b1), .IN2(~na184_1), .IN3(1'b1), .IN4(~na196_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x39y89     80'h00_FE00_00_0000_0CEE_D000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a224_1 ( .OUT(na224_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na44_1), .IN8(na1345_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a224_2 ( .OUT(na224_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na224_1_i) );
// C_MX2b////      x39y88     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a225_1 ( .OUT(na225_1), .IN1(1'b1), .IN2(~na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1346_2), .IN8(~na826_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x31y92     80'h00_0018_00_0040_0C0A_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a226_1 ( .OUT(na226_1), .IN1(1'b0), .IN2(na160_1), .IN3(1'b0), .IN4(na1347_2), .IN5(~na166_1), .IN6(1'b1), .IN7(~na167_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x35y102     80'h00_FE00_80_0000_0C88_ACAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a227_1 ( .OUT(na227_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1348_1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a227_2 ( .OUT(na227_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na227_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a227_4 ( .OUT(na227_2_i), .IN1(na1558_2), .IN2(1'b1), .IN3(na1313_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a227_5 ( .OUT(na227_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na227_2_i) );
// C_MX2b////      x32y100     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a228_1 ( .OUT(na228_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1615_2), .IN5(~na1349_2), .IN6(1'b0), .IN7(~na818_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x37y86     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a229_4 ( .OUT(na229_2_i), .IN1(na1350_1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a229_5 ( .OUT(na229_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na229_2_i) );
// C_MX2b////      x33y87     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a230_1 ( .OUT(na230_1), .IN1(1'b1), .IN2(~na256_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1351_1), .IN6(na229_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x27y107     80'h00_FE00_80_0000_0C88_A5A3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a231_1 ( .OUT(na231_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na232_1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a231_2 ( .OUT(na231_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na231_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a231_4 ( .OUT(na231_2_i), .IN1(1'b1), .IN2(~na304_1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a231_5 ( .OUT(na231_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na231_2_i) );
// C_MX2b////      x25y109     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a232_1 ( .OUT(na232_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1610_2), .IN5(~na231_1), .IN6(1'b0), .IN7(~na1352_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x31y110     80'h00_0018_00_0000_0888_88CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a233_1 ( .OUT(na233_1), .IN1(na237_1), .IN2(1'b1), .IN3(1'b1), .IN4(na300_2), .IN5(na299_2), .IN6(na234_1), .IN7(na1627_2),
                     .IN8(na300_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x31y106     80'h00_0018_00_0000_0C88_38FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a234_1 ( .OUT(na234_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1363_2), .IN6(na371_1), .IN7(1'b1), .IN8(~na292_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x25y116     80'h00_0018_00_0000_0888_8882
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a235_1 ( .OUT(na235_1), .IN1(na299_2), .IN2(~na1624_2), .IN3(na1627_2), .IN4(na300_1), .IN5(na297_2), .IN6(na293_2), .IN7(na298_1),
                     .IN8(na300_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x27y115     80'h00_0018_00_0000_0C88_28FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a237_1 ( .OUT(na237_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na297_2), .IN6(na293_2), .IN7(na298_1), .IN8(~na1625_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x23y107     80'h00_0018_00_0000_0888_8848
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a238_1 ( .OUT(na238_1), .IN1(na231_1), .IN2(na316_1), .IN3(~na314_1), .IN4(na318_1), .IN5(na231_2), .IN6(na316_2), .IN7(na314_2),
                     .IN8(na318_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x32y105     80'h00_FE00_00_0000_0CEE_D000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a241_1 ( .OUT(na241_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na44_1), .IN8(na1353_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a241_2 ( .OUT(na241_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na241_1_i) );
// C_///ORAND/      x32y110     80'h00_0060_00_0000_0C08_FFBB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a242_4 ( .OUT(na242_2), .IN1(na23_1), .IN2(~na1152_1), .IN3(na241_1), .IN4(~na36_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x21y85     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a244_4 ( .OUT(na244_2_i), .IN1(na1357_1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a244_5 ( .OUT(na244_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na244_2_i) );
// C_AND////      x28y107     80'h00_0018_00_0000_0C88_14FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a246_1 ( .OUT(na246_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na23_1), .IN6(na1621_2), .IN7(~na276_1), .IN8(~na1_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x19y98     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a247_1 ( .OUT(na247_1), .IN1(1'b1), .IN2(~na1359_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1706_2), .IN8(~na335_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y102     80'h00_0060_00_0000_0C08_FF84
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a248_4 ( .OUT(na248_2), .IN1(~na23_1), .IN2(na173_2), .IN3(na1622_2), .IN4(na1_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x27y103     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a249_1 ( .OUT(na249_1), .IN1(1'b1), .IN2(na1621_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1153_1), .IN6(~na1360_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x30y101     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a250_4 ( .OUT(na250_2), .IN1(na23_1), .IN2(1'b1), .IN3(na241_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x30y107     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a251_1 ( .OUT(na251_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na297_1), .IN6(1'b0), .IN7(na314_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x30y110     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a252_4 ( .OUT(na252_2), .IN1(1'b1), .IN2(na293_2), .IN3(na251_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y102     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a253_1 ( .OUT(na253_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1582_2), .IN8(na1_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x23y99     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a254_4 ( .OUT(na254_2_i), .IN1(na1361_1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a254_5 ( .OUT(na254_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na254_2_i) );
// C_MX2b////      x23y104     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a255_1 ( .OUT(na255_1), .IN1(1'b1), .IN2(na1359_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na359_2), .IN6(~na1154_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x33y94     80'h00_FE00_00_0000_0888_FEA5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a256_1 ( .OUT(na256_1_i), .IN1(~na257_1), .IN2(1'b0), .IN3(na44_1), .IN4(1'b0), .IN5(na1691_2), .IN6(na256_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a256_2 ( .OUT(na256_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na256_1_i) );
// C_AND////      x25y103     80'h00_0018_00_0000_0888_3584
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a257_1 ( .OUT(na257_1), .IN1(~na1363_1), .IN2(na1707_2), .IN3(na276_1), .IN4(na292_1), .IN5(~na23_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na1_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x25y95     80'h00_FE00_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a258_1 ( .OUT(na258_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na44_1), .IN8(~na259_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a258_2 ( .OUT(na258_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na258_1_i) );
// C_MX2b////      x24y94     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a259_1 ( .OUT(na259_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1561_2), .IN5(~na258_1), .IN6(1'b0), .IN7(~na772_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x25y96     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a260_1 ( .OUT(na260_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1364_1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a260_2 ( .OUT(na260_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na260_1_i) );
// C_AND///AND/      x29y99     80'h00_0078_00_0000_0C88_CC5A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a262_1 ( .OUT(na262_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1621_2), .IN7(1'b1), .IN8(na1365_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a262_4 ( .OUT(na262_2), .IN1(na1363_2), .IN2(1'b1), .IN3(~na246_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x38y97     80'h00_FE00_80_0000_0C88_AC8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a263_1 ( .OUT(na263_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1366_1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a263_2 ( .OUT(na263_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na263_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a263_4 ( .OUT(na263_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na44_1), .IN4(na1378_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a263_5 ( .OUT(na263_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na263_2_i) );
// C_MX2b////      x34y100     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a264_1 ( .OUT(na264_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1615_2), .IN5(1'b0), .IN6(~na1367_1), .IN7(1'b0), .IN8(~na816_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x43y109     80'h00_FE00_00_0000_0888_FE5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a265_1 ( .OUT(na265_1_i), .IN1(1'b0), .IN2(na470_2), .IN3(~na266_1), .IN4(1'b0), .IN5(na265_1), .IN6(na1671_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a265_2 ( .OUT(na265_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na265_1_i) );
// C_AND////      x44y103     80'h00_0018_00_0000_0888_43F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a266_1 ( .OUT(na266_1), .IN1(na397_2), .IN2(na267_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na267_2), .IN7(~na25_1),
                     .IN8(na13_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x43y104     80'h00_0078_00_0000_0C88_CCC3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a267_1 ( .OUT(na267_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1441_2), .IN7(1'b1), .IN8(na13_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a267_4 ( .OUT(na267_2), .IN1(1'b1), .IN2(~na269_1), .IN3(1'b1), .IN4(na1143_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x45y116     80'h00_0018_00_0040_0CE9_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a269_1 ( .OUT(na269_1), .IN1(na1371_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1370_1), .IN5(~na1141_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na1138_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x36y108     80'h00_FE00_80_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a270_1 ( .OUT(na270_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1372_1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a270_2 ( .OUT(na270_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na270_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a270_4 ( .OUT(na270_2_i), .IN1(1'b1), .IN2(na1383_1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a270_5 ( .OUT(na270_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na270_2_i) );
// C_ORAND////      x36y113     80'h00_0018_00_0000_0C88_7BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a271_1 ( .OUT(na271_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na23_1), .IN6(~na1155_1), .IN7(~na1679_2), .IN8(~na36_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x38y103     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a272_4 ( .OUT(na272_2_i), .IN1(na1375_1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a272_5 ( .OUT(na272_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na272_2_i) );
// C_///ORAND/      x38y114     80'h00_0060_00_0000_0C08_FF7B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a273_4 ( .OUT(na273_2), .IN1(na23_1), .IN2(~na1156_1), .IN3(~na1677_2), .IN4(~na36_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y97     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a275_1 ( .OUT(na275_1), .IN1(1'b1), .IN2(~na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1379_1), .IN8(~na816_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x30y101     80'h00_FE00_00_0000_0C88_ADFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a276_1 ( .OUT(na276_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1380_2), .IN6(na1381_2), .IN7(na44_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a276_2 ( .OUT(na276_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na276_1_i) );
// C_ORAND////      x36y107     80'h00_0018_00_0000_0C88_7BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a281_1 ( .OUT(na281_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na23_1), .IN6(~na1157_1), .IN7(~na1676_2), .IN8(~na36_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x52y103     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a282_4 ( .OUT(na282_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(na1386_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a282_5 ( .OUT(na282_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na282_2_i) );
// C_MX2b////      x54y112     80'h00_0018_00_0040_0AC4_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a283_1 ( .OUT(na283_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na717_2), .IN8(na284_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x52y116     80'h00_0018_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_1 ( .OUT(na284_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na286_2), .IN7(~na1387_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x49y116     80'h00_0060_00_0000_0C08_FF48
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a286_4 ( .OUT(na286_2), .IN1(na1141_1), .IN2(na1136_1), .IN3(~na1701_2), .IN4(na1138_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x49y98     80'h00_FE00_00_0000_0CEE_0B00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a287_1 ( .OUT(na287_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1388_1), .IN6(~na470_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a287_2 ( .OUT(na287_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na287_1_i) );
// C_ORAND///ORAND/      x49y104     80'h00_0078_00_0000_0C88_3B3D
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a288_1 ( .OUT(na288_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na265_1), .IN6(~na1669_2), .IN7(1'b0), .IN8(~na289_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a288_4 ( .OUT(na288_2), .IN1(~na265_1), .IN2(na1234_1), .IN3(1'b0), .IN4(~na70_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x52y116     80'h00_0060_00_0000_0C08_FF4C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a289_4 ( .OUT(na289_2), .IN1(1'b1), .IN2(na1136_1), .IN3(~na1246_1), .IN4(na290_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x52y114     80'h00_0018_00_0000_0C88_38FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a290_1 ( .OUT(na290_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(na1616_2), .IN7(1'b1), .IN8(~na1143_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND*/D      x23y117     80'h00_FE00_80_0000_0C07_FF55
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a291_4 ( .OUT(na291_2_i), .IN1(~na291_2), .IN2(1'b1), .IN3(~na752_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a291_5 ( .OUT(na291_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na291_2_i) );
// C_ORAND*/D///      x30y102     80'h00_FE00_00_0000_0388_ABFF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a292_1 ( .OUT(na292_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na56_1), .IN6(~na1621_2), .IN7(na44_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a292_2 ( .OUT(na292_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na292_1_i) );
// C_///ORAND*/D      x29y112     80'h00_FE00_80_0000_0C07_FF77
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a293_4 ( .OUT(na293_2_i), .IN1(~na1623_2), .IN2(~na294_2), .IN3(~na295_1), .IN4(~na1685_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a293_5 ( .OUT(na293_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na293_2_i) );
// C_///AND/      x29y110     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a294_4 ( .OUT(na294_2), .IN1(1'b1), .IN2(~na234_1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x30y109     80'h00_0018_00_0000_0C88_A2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a295_1 ( .OUT(na295_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1611_2), .IN6(~na235_1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D//ORAND*/D      x29y111     80'h00_FE00_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a297_1 ( .OUT(na297_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na297_1), .IN6(~na294_2), .IN7(~na295_1),
                     .IN8(~na1684_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a297_2 ( .OUT(na297_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na297_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a297_4 ( .OUT(na297_2_i), .IN1(~na297_2), .IN2(~na294_2), .IN3(~na295_1), .IN4(~na798_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a297_5 ( .OUT(na297_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na297_2_i) );
// C_ORAND*/D///      x24y113     80'h00_FE00_00_0000_0388_77FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a298_1 ( .OUT(na298_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1626_2), .IN6(~na294_2), .IN7(~na295_1),
                     .IN8(~na798_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a298_2 ( .OUT(na298_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na298_1_i) );
// C_ORAND*/D//ORAND*/D      x25y113     80'h00_FE00_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a299_1 ( .OUT(na299_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na299_1), .IN6(~na294_2), .IN7(~na295_1),
                     .IN8(~na1683_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a299_2 ( .OUT(na299_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na299_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a299_4 ( .OUT(na299_2_i), .IN1(~na299_2), .IN2(~na294_2), .IN3(~na295_1), .IN4(~na794_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a299_5 ( .OUT(na299_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na299_2_i) );
// C_ORAND*/D//ORAND*/D      x28y116     80'h00_FE00_80_0000_0387_77D7
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a300_1 ( .OUT(na300_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1628_2), .IN6(~na294_2), .IN7(~na295_1),
                     .IN8(~na794_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a300_2 ( .OUT(na300_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na300_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a300_4 ( .OUT(na300_2_i), .IN1(~na1629_2), .IN2(~na294_2), .IN3(~na295_1), .IN4(na300_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a300_5 ( .OUT(na300_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na300_2_i) );
// C_MX2b////      x25y110     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a304_1 ( .OUT(na304_1), .IN1(1'b1), .IN2(na233_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na231_2), .IN6(~na1408_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x25y108     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a306_1 ( .OUT(na306_1), .IN1(1'b1), .IN2(~na233_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1409_2), .IN6(~na316_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x25y107     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a308_1 ( .OUT(na308_1), .IN1(1'b1), .IN2(~na233_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1410_1), .IN8(~na318_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x50y90     80'h00_FE00_80_0000_0C88_ACCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a309_1 ( .OUT(na309_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1411_1), .IN7(na1650_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a309_2 ( .OUT(na309_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na309_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a309_4 ( .OUT(na309_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(1'b1), .IN4(na1439_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a309_5 ( .OUT(na309_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na309_2_i) );
// C_AND///AND/      x51y85     80'h00_0078_00_0000_0C88_5CAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a311_1 ( .OUT(na311_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na701_1), .IN7(~na312_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a311_4 ( .OUT(na311_2), .IN1(1'b1), .IN2(na48_2), .IN3(na49_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x52y87     80'h00_0018_00_0000_0888_8AC8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a312_1 ( .OUT(na312_1), .IN1(na353_1), .IN2(na355_2), .IN3(1'b1), .IN4(na309_2), .IN5(na353_2), .IN6(1'b1), .IN7(na324_2),
                     .IN8(na309_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x32y107     80'h00_FE00_80_0000_0C88_2FA3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a314_1 ( .OUT(na314_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na44_1), .IN8(~na315_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a314_2 ( .OUT(na314_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na314_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a314_4 ( .OUT(na314_2_i), .IN1(1'b1), .IN2(~na321_1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a314_5 ( .OUT(na314_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na314_2_i) );
// C_MX2b////      x28y108     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a315_1 ( .OUT(na315_1), .IN1(1'b1), .IN2(na233_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na314_1), .IN8(~na1412_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x25y106     80'h00_FE00_80_0000_0C88_2FA3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a316_1 ( .OUT(na316_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na44_1), .IN8(~na317_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a316_2 ( .OUT(na316_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na316_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a316_4 ( .OUT(na316_2_i), .IN1(1'b1), .IN2(~na306_1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a316_5 ( .OUT(na316_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na316_2_i) );
// C_MX2b////      x24y108     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a317_1 ( .OUT(na317_1), .IN1(1'b1), .IN2(~na233_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1413_2), .IN6(~na316_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x28y106     80'h00_FE00_80_0000_0C88_5AA5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a318_1 ( .OUT(na318_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1558_2), .IN6(1'b1), .IN7(~na319_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a318_2 ( .OUT(na318_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na318_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a318_4 ( .OUT(na318_2_i), .IN1(~na308_1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a318_5 ( .OUT(na318_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na318_2_i) );
// C_MX2b////      x24y107     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a319_1 ( .OUT(na319_1), .IN1(1'b1), .IN2(~na233_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1414_1), .IN8(~na318_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x29y108     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a321_1 ( .OUT(na321_1), .IN1(1'b1), .IN2(na233_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na314_2), .IN8(~na1415_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x24y95     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a322_1 ( .OUT(na322_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na44_1), .IN8(na1416_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a322_2 ( .OUT(na322_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na322_1_i) );
// C_AND/D//AND/D      x24y96     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a323_1 ( .OUT(na323_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1417_1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a323_2 ( .OUT(na323_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na323_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a323_4 ( .OUT(na323_2_i), .IN1(na1356_1), .IN2(1'b1), .IN3(na44_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a323_5 ( .OUT(na323_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na323_2_i) );
// C_///AND/D      x52y95     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a324_4 ( .OUT(na324_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(na1418_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a324_5 ( .OUT(na324_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na324_2_i) );
// C_AND////      x52y96     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a325_1 ( .OUT(na325_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na699_2), .IN6(1'b1), .IN7(~na312_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/D      x23y95     80'h00_FE00_80_0000_0C08_FFA6
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a328_4 ( .OUT(na328_2_i), .IN1(na328_2), .IN2(~na57_2), .IN3(~na44_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a328_5 ( .OUT(na328_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na328_2_i) );
// C_///AND/      x46y85     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a330_4 ( .OUT(na330_2), .IN1(na703_1), .IN2(1'b1), .IN3(~na49_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP/D///      x48y97     80'h00_FE00_00_0000_0C88_6CFF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a331_1 ( .OUT(na331_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na470_2), .IN7(na331_1), .IN8(~na13_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a331_2 ( .OUT(na331_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na331_1_i) );
// C_///AND/      x27y105     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a332_4 ( .OUT(na332_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na251_1), .IN4(na318_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y106     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a333_4 ( .OUT(na333_2), .IN1(na299_1), .IN2(1'b1), .IN3(na251_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x30y99     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a334_1 ( .OUT(na334_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na171_1), .IN7(1'b1), .IN8(na1_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x22y98     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a335_1 ( .OUT(na335_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1424_1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a335_2 ( .OUT(na335_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na335_1_i) );
// C_MX2b////      x24y101     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a336_1 ( .OUT(na336_1), .IN1(1'b1), .IN2(na1359_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na341_1), .IN6(~na1158_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x47y88     80'h00_FE00_80_0000_0C88_F8A4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a337_1 ( .OUT(na337_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1425_1), .IN6(na470_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a337_2 ( .OUT(na337_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na337_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a337_4 ( .OUT(na337_2_i), .IN1(~na311_2), .IN2(na470_2), .IN3(na1419_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a337_5 ( .OUT(na337_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na337_2_i) );
// C_///AND/      x39y89     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a338_4 ( .OUT(na338_2), .IN1(1'b1), .IN2(na705_2), .IN3(~na49_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x27y106     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a339_1 ( .OUT(na339_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na316_2), .IN7(~na251_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x26y100     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a340_4 ( .OUT(na340_2), .IN1(na170_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x23y97     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a341_1 ( .OUT(na341_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na44_1), .IN8(na1426_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a341_2 ( .OUT(na341_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na341_1_i) );
// C_MX2b////      x31y102     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a342_1 ( .OUT(na342_1), .IN1(1'b1), .IN2(na1359_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na347_1), .IN6(~na1159_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x42y88     80'h00_FE00_80_0000_0C88_ACCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a343_1 ( .OUT(na343_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(na1427_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a343_2 ( .OUT(na343_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na343_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a343_4 ( .OUT(na343_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(1'b1), .IN4(na1422_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a343_5 ( .OUT(na343_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na343_2_i) );
// C_///AND/      x46y93     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a344_4 ( .OUT(na344_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na49_1), .IN4(~na343_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y107     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a345_1 ( .OUT(na345_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na297_1), .IN6(1'b1), .IN7(na314_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x34y103     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a346_4 ( .OUT(na346_2), .IN1(1'b1), .IN2(1'b1), .IN3(na167_1), .IN4(na1_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x23y99     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a347_1 ( .OUT(na347_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1428_1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a347_2 ( .OUT(na347_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na347_1_i) );
// C_MX2b////      x26y103     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a348_1 ( .OUT(na348_1), .IN1(1'b1), .IN2(na1359_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na351_1), .IN6(~na1160_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x26y104     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a349_1 ( .OUT(na349_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na316_1), .IN7(~na251_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x31y104     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a350_4 ( .OUT(na350_2), .IN1(na166_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x25y99     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a351_1 ( .OUT(na351_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1429_1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a351_2 ( .OUT(na351_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na351_1_i) );
// C_MX2b////      x23y102     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a352_1 ( .OUT(na352_1), .IN1(1'b1), .IN2(na1359_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na254_2), .IN6(~na1161_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x49y89     80'h00_FE00_80_0000_0C88_F8AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a353_1 ( .OUT(na353_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1430_1), .IN6(na470_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a353_2 ( .OUT(na353_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na353_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a353_4 ( .OUT(na353_2_i), .IN1(1'b1), .IN2(na1433_1), .IN3(na1650_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a353_5 ( .OUT(na353_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na353_2_i) );
// C_AND////      x51y94     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a354_1 ( .OUT(na354_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na699_1), .IN6(1'b1), .IN7(~na312_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x53y96     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a355_4 ( .OUT(na355_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(na1431_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a355_5 ( .OUT(na355_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na355_2_i) );
// C_///AND/      x51y87     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a356_4 ( .OUT(na356_2), .IN1(1'b1), .IN2(na697_2), .IN3(~na312_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y106     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a357_1 ( .OUT(na357_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na297_2), .IN6(1'b1), .IN7(na251_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x34y102     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a358_4 ( .OUT(na358_2), .IN1(1'b1), .IN2(na160_1), .IN3(1'b1), .IN4(na1_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x25y99     80'h00_FE00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a359_4 ( .OUT(na359_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na44_1), .IN4(na1432_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a359_5 ( .OUT(na359_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na359_2_i) );
// C_MX2b////      x28y103     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a360_1 ( .OUT(na360_1), .IN1(1'b1), .IN2(~na1359_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1162_1), .IN8(~na365_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x51y88     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a362_1 ( .OUT(na362_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na697_1), .IN7(~na312_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y105     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a363_4 ( .OUT(na363_2), .IN1(na1614_2), .IN2(1'b1), .IN3(na298_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y99     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a364_1 ( .OUT(na364_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na167_2), .IN8(na1_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x22y98     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a365_4 ( .OUT(na365_2_i), .IN1(na1558_2), .IN2(1'b1), .IN3(na1434_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a365_5 ( .OUT(na365_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na365_2_i) );
// C_AND///AND/      x21y98     80'h00_0078_00_0000_0C88_CC54
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a366_1 ( .OUT(na366_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1359_2), .IN7(1'b1), .IN8(na1163_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a366_4 ( .OUT(na366_2), .IN1(~na328_2), .IN2(na57_2), .IN3(~na1358_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x44y96     80'h00_FE00_80_0000_0C88_CCF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a367_1 ( .OUT(na367_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1), .IN8(na1435_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a367_2 ( .OUT(na367_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na367_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a367_4 ( .OUT(na367_2_i), .IN1(na1531_1), .IN2(na470_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a367_5 ( .OUT(na367_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na367_2_i) );
// C_OR/D///      x22y87     80'h00_FE00_00_0000_0CEE_5C00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a368_1 ( .OUT(na368_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1436_1), .IN7(~na44_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a368_2 ( .OUT(na368_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na368_1_i) );
// C_///ORAND/      x27y100     80'h00_0060_00_0000_0C08_FFC7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a369_4 ( .OUT(na369_2), .IN1(~na39_2), .IN2(~na1382_1), .IN3(1'b0), .IN4(na1708_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x30y100     80'h00_0018_00_0000_0C88_4AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a370_1 ( .OUT(na370_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na23_1), .IN6(1'b1), .IN7(~na241_1), .IN8(na292_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x29y104     80'h00_FE00_00_0040_0C03_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a371_1 ( .OUT(na371_1_i), .IN1(na1437_1), .IN2(na371_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1621_2), .IN7(~na44_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a371_2 ( .OUT(na371_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na371_1_i) );
// C_AND/D///      x47y93     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a372_1 ( .OUT(na372_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(na1438_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a372_2 ( .OUT(na372_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na372_1_i) );
// C_///AND/      x52y93     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a374_4 ( .OUT(na374_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na312_1), .IN4(~na309_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x24y91     80'h00_FE18_00_0000_0888_AFF5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a375_1 ( .OUT(na375_1), .IN1(~na376_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a375_5 ( .OUT(na375_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na375_1) );
// C_MX2b////      x21y89     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a376_1 ( .OUT(na376_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na375_2), .IN8(~na770_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x23y92     80'h00_FE18_00_0000_0888_AFF5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a377_1 ( .OUT(na377_1), .IN1(~na378_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na44_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a377_5 ( .OUT(na377_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na377_1) );
// C_MX2b////      x23y91     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a378_1 ( .OUT(na378_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1561_2), .IN5(1'b0), .IN6(~na377_2), .IN7(1'b0), .IN8(~na770_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x50y91     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a379_4 ( .OUT(na379_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(na1440_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a379_5 ( .OUT(na379_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na379_2_i) );
// C_MX2b////      x50y92     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a380_1 ( .OUT(na380_1), .IN1(1'b1), .IN2(na1441_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na451_1), .IN6(na1441_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x43y99     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a381_1 ( .OUT(na381_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1147_1), .IN6(1'b1), .IN7(na25_1), .IN8(na13_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x46y92     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a382_1 ( .OUT(na382_1), .IN1(1'b1), .IN2(na1646_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1164_1), .IN8(~na1442_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x45y93     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a383_1 ( .OUT(na383_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na32_1), .IN7(1'b1), .IN8(na416_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x49y96     80'h00_0018_00_0000_0888_F7C3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a384_1 ( .OUT(na384_1), .IN1(1'b0), .IN2(~na1632_2), .IN3(1'b0), .IN4(na13_1), .IN5(~na69_2), .IN6(~na1441_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x51y97     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a385_4 ( .OUT(na385_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(na1444_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a385_5 ( .OUT(na385_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na385_2_i) );
// C_MX2b////      x49y106     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a386_1 ( .OUT(na386_1), .IN1(~na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1445_2), .IN8(~na730_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x51y118     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a388_4 ( .OUT(na388_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(na1447_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a388_5 ( .OUT(na388_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na388_2_i) );
// C_///AND/      x45y108     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a389_4 ( .OUT(na389_2), .IN1(~na69_2), .IN2(na267_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x43y97     80'h00_0018_00_0000_0CEE_3A00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a390_1 ( .OUT(na390_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1448_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na420_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x47y97     80'h00_FE00_80_0000_0C88_ACF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a391_1 ( .OUT(na391_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(na1449_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a391_2 ( .OUT(na391_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na391_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a391_4 ( .OUT(na391_2_i), .IN1(na1451_1), .IN2(na470_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a391_5 ( .OUT(na391_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na391_2_i) );
// C_MX2b////      x47y104     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a392_1 ( .OUT(na392_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na720_2), .IN8(~na1450_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y106     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a394_1 ( .OUT(na394_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na720_1), .IN8(~na1452_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x45y118     80'h00_0018_00_0000_0C88_21FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a395_1 ( .OUT(na395_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1141_1), .IN6(~na1136_1), .IN7(na1133_1),
                     .IN8(~na1138_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x52y115     80'h00_FE00_00_0000_0C88_ECFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a396_1 ( .OUT(na396_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na470_2), .IN7(na396_1), .IN8(na13_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a396_2 ( .OUT(na396_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na396_1_i) );
// C_///ORAND*/D      x45y101     80'h00_FE00_80_0000_0C07_FF37
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a397_4 ( .OUT(na397_2_i), .IN1(~na1150_1), .IN2(~na400_2), .IN3(1'b0), .IN4(~na1455_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a397_5 ( .OUT(na397_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na397_2_i) );
// C_///AND/      x41y100     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a399_4 ( .OUT(na399_2), .IN1(1'b1), .IN2(na1441_2), .IN3(na1647_2), .IN4(na13_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x39y108     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a400_4 ( .OUT(na400_2), .IN1(na383_1), .IN2(na267_1), .IN3(na1651_2), .IN4(na420_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x39y95     80'h00_FE00_80_0000_0C88_F8AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a402_1 ( .OUT(na402_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1457_1), .IN6(na470_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a402_2 ( .OUT(na402_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na402_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a402_4 ( .OUT(na402_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(na1469_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a402_5 ( .OUT(na402_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na402_2_i) );
// C_ORAND////      x40y99     80'h00_0018_00_0000_0C88_7DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a403_1 ( .OUT(na403_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1165_1), .IN6(na32_1), .IN7(~na404_1), .IN8(~na1666_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x42y95     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a404_1 ( .OUT(na404_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na32_1), .IN7(~na405_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x42y113     80'h00_0018_00_0000_0888_1154
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a405_1 ( .OUT(na405_1), .IN1(~na1147_1), .IN2(na407_2), .IN3(~na1697_2), .IN4(1'b1), .IN5(~na1141_1), .IN6(~na1700_2), .IN7(~na1133_1),
                     .IN8(~na1138_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x41y114     80'h00_0060_00_0000_0C08_FFC1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a407_4 ( .OUT(na407_2), .IN1(~na1150_1), .IN2(~na1146_1), .IN3(1'b1), .IN4(na416_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x39y100     80'h00_0060_00_0000_0C08_FF7D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a409_4 ( .OUT(na409_2), .IN1(~na1166_1), .IN2(na32_1), .IN3(~na404_1), .IN4(~na1662_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x37y104     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a410_1 ( .OUT(na410_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1), .IN8(na1463_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a410_2 ( .OUT(na410_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na410_1_i) );
// C_ORAND////      x41y99     80'h00_0018_00_0000_0C88_7DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a411_1 ( .OUT(na411_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1167_1), .IN6(na32_1), .IN7(~na404_1), .IN8(~na1664_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x39y101     80'h00_FE00_80_0000_0C88_F8AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a412_1 ( .OUT(na412_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1466_1), .IN6(na470_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a412_2 ( .OUT(na412_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na412_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a412_4 ( .OUT(na412_2_i), .IN1(1'b1), .IN2(na1460_1), .IN3(na1650_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a412_5 ( .OUT(na412_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na412_2_i) );
// C_///ORAND/      x39y102     80'h00_0060_00_0000_0C08_FF7D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a413_4 ( .OUT(na413_2), .IN1(~na1168_1), .IN2(na32_1), .IN3(~na404_1), .IN4(~na1663_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x42y97     80'h00_0018_00_0000_0C88_7DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a415_1 ( .OUT(na415_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1169_1), .IN6(na32_1), .IN7(~na404_1), .IN8(~na1660_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x46y98     80'h00_FE00_00_0000_0CEE_C300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a416_1 ( .OUT(na416_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na470_2), .IN7(1'b0), .IN8(na1472_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a416_2 ( .OUT(na416_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na416_1_i) );
// C_///ORAND/      x44y99     80'h00_0060_00_0000_0C08_FFDD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a417_4 ( .OUT(na417_2), .IN1(~na1170_1), .IN2(na32_1), .IN3(~na404_1), .IN4(na416_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x46y98     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a418_4 ( .OUT(na418_2_i), .IN1(na1475_1), .IN2(na470_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a418_5 ( .OUT(na418_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na418_2_i) );
// C_MX2b////      x42y105     80'h00_0018_00_0040_0AC4_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a419_1 ( .OUT(na419_1), .IN1(~na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1476_1), .IN8(na418_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND*/D      x42y96     80'h00_FE00_80_0000_0C07_FFBC
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a420_4 ( .OUT(na420_2_i), .IN1(1'b0), .IN2(na470_2), .IN3(na1478_2), .IN4(~na420_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a420_5 ( .OUT(na420_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na420_2_i) );
// C_AND/D//AND/D      x46y110     80'h00_FE00_80_0000_0C88_ACF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a421_1 ( .OUT(na421_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1479_1), .IN7(na1650_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a421_2 ( .OUT(na421_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na421_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a421_4 ( .OUT(na421_2_i), .IN1(na1482_1), .IN2(na470_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a421_5 ( .OUT(na421_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na421_2_i) );
// C_MX2b////      x46y111     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a422_1 ( .OUT(na422_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na726_2), .IN8(~na1480_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y111     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a425_1 ( .OUT(na425_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na726_1), .IN8(~na1483_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x49y118     80'h00_0018_00_0040_0CF9_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a426_1 ( .OUT(na426_1), .IN1(~na1371_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1484_2), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na1138_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x52y108     80'h00_FE00_80_0000_0C88_ACF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a427_1 ( .OUT(na427_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(na1486_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a427_2 ( .OUT(na427_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na427_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a427_4 ( .OUT(na427_2_i), .IN1(na1489_1), .IN2(na470_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a427_5 ( .OUT(na427_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na427_2_i) );
// C_MX2b////      x52y111     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a428_1 ( .OUT(na428_1), .IN1(~na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1487_1), .IN8(~na724_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x49y117     80'h00_0018_00_0040_0CFC_5500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a429_1 ( .OUT(na429_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1274_2), .IN4(~na1138_1), .IN5(~na1141_1), .IN6(1'b1), .IN7(~na1697_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y113     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a431_1 ( .OUT(na431_1), .IN1(~na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1490_1), .IN8(~na724_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x46y105     80'h00_FE00_80_0000_0C88_CCAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a432_1 ( .OUT(na432_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1), .IN8(na1491_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a432_2 ( .OUT(na432_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na432_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a432_4 ( .OUT(na432_2_i), .IN1(1'b1), .IN2(na1493_1), .IN3(na1650_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a432_5 ( .OUT(na432_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na432_2_i) );
// C_MX2b////      x46y112     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a433_1 ( .OUT(na433_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na722_2), .IN8(~na1492_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x46y114     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a435_1 ( .OUT(na435_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na722_1), .IN8(~na1494_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x45y104     80'h00_FE00_80_0000_0C88_F8CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a436_1 ( .OUT(na436_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1495_1), .IN6(na470_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a436_2 ( .OUT(na436_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na436_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a436_4 ( .OUT(na436_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(1'b1), .IN4(na1497_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a436_5 ( .OUT(na436_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na436_2_i) );
// C_MX2b////      x47y109     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a437_1 ( .OUT(na437_1), .IN1(~na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1496_1), .IN8(~na719_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x45y111     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a439_1 ( .OUT(na439_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1498_1), .IN6(na440_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x43y112     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a440_1 ( .OUT(na440_1), .IN1(~na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1500_1), .IN8(~na719_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/D      x51y102     80'h00_FE00_80_0000_0C0E_FFA3
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a441_4 ( .OUT(na441_2_i), .IN1(1'b0), .IN2(~na470_2), .IN3(na1501_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a441_5 ( .OUT(na441_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na441_2_i) );
// C_MX2b////      x49y111     80'h00_0018_00_0040_0AC4_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a442_1 ( .OUT(na442_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na717_1), .IN8(na443_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y118     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a443_1 ( .OUT(na443_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1143_1), .IN5(1'b0), .IN6(~na395_1), .IN7(1'b0), .IN8(~na1502_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x43y111     80'h00_0018_00_0000_0C88_7BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a446_1 ( .OUT(na446_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na265_1), .IN6(~na1670_2), .IN7(~na1506_1),
                     .IN8(~na290_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x47y90     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a448_4 ( .OUT(na448_2), .IN1(1'b0), .IN2(na337_1), .IN3(na324_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x45y91     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a449_1 ( .OUT(na449_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na353_1), .IN6(~na448_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x42y103     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a450_4 ( .OUT(na450_2), .IN1(1'b1), .IN2(na1146_1), .IN3(na25_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x49y93     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a451_1 ( .OUT(na451_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1507_1), .IN6(na470_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a451_2 ( .OUT(na451_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na451_1_i) );
// C_MX2b////      x47y92     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a452_1 ( .OUT(na452_1), .IN1(1'b1), .IN2(na1441_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na489_2), .IN6(~na1171_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x43y110     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a453_4 ( .OUT(na453_2_i), .IN1(na1508_1), .IN2(na470_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a453_5 ( .OUT(na453_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na453_2_i) );
// C_///ORAND/      x51y113     80'h00_0060_00_0000_0C08_FF7B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a454_4 ( .OUT(na454_2), .IN1(na265_1), .IN2(~na1668_2), .IN3(~na1510_1), .IN4(~na290_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x51y103     80'h00_FE00_00_0000_0CEE_C300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a456_1 ( .OUT(na456_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na470_2), .IN7(1'b0), .IN8(na1511_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a456_2 ( .OUT(na456_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na456_1_i) );
// C_///ORAND/      x51y112     80'h00_0060_00_0000_0C08_FF3B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a457_4 ( .OUT(na457_2), .IN1(na265_1), .IN2(~na1667_2), .IN3(1'b0), .IN4(~na458_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x54y116     80'h00_0060_00_0000_0C08_FF43
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a458_4 ( .OUT(na458_2), .IN1(1'b1), .IN2(~na1136_1), .IN3(~na1246_1), .IN4(na290_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x49y97     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a459_4 ( .OUT(na459_2_i), .IN1(1'b1), .IN2(na1514_1), .IN3(na1650_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a459_5 ( .OUT(na459_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na459_2_i) );
// C_MX2b////      x47y108     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a460_1 ( .OUT(na460_1), .IN1(~na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1515_1), .IN8(~na711_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x51y100     80'h00_FE00_80_0000_0C88_CCF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a461_1 ( .OUT(na461_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1), .IN8(na1516_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a461_2 ( .OUT(na461_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na461_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a461_4 ( .OUT(na461_2_i), .IN1(na1518_1), .IN2(na470_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a461_5 ( .OUT(na461_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na461_2_i) );
// C_MX2b////      x47y113     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a462_1 ( .OUT(na462_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na736_2), .IN8(~na1517_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y107     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a464_1 ( .OUT(na464_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na736_1), .IN8(~na1519_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x51y97     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a465_1 ( .OUT(na465_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(na1520_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a465_2 ( .OUT(na465_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na465_1_i) );
// C_MX2b////      x49y108     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a466_1 ( .OUT(na466_1), .IN1(~na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1521_1), .IN8(~na734_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x47y89     80'h00_FE00_00_0040_0C05_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a467_1 ( .OUT(na467_1_i), .IN1(na467_1), .IN2(1'b0), .IN3(na1522_2), .IN4(1'b0), .IN5(1'b1), .IN6(~na470_2), .IN7(1'b1),
                     .IN8(~na420_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a467_2 ( .OUT(na467_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na467_1_i) );
// C_ORAND*/D///      x52y107     80'h00_FE00_00_0000_0788_FCDD
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a468_1 ( .OUT(na468_1_i), .IN1(~na1562_2), .IN2(na470_1), .IN3(~na468_1), .IN4(na1524_1), .IN5(1'b0), .IN6(na470_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a468_2 ( .OUT(na468_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na468_1_i) );
// C_AND///AND/      x43y98     80'h00_0078_00_0000_0C88_CC5A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a470_1 ( .OUT(na470_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na32_1), .IN7(1'b1), .IN8(na420_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a470_4 ( .OUT(na470_2), .IN1(na1178_1), .IN2(1'b1), .IN3(~na529_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x47y90     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a471_1 ( .OUT(na471_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na337_1), .IN7(~na324_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x44y108     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a472_4 ( .OUT(na472_2), .IN1(1'b1), .IN2(1'b1), .IN3(na25_1), .IN4(na1696_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x46y90     80'h00_FE00_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a473_4 ( .OUT(na473_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(1'b1), .IN4(~na474_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a473_5 ( .OUT(na473_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na473_2_i) );
// C_MX2b////      x50y96     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a474_1 ( .OUT(na474_1), .IN1(1'b1), .IN2(~na384_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1525_2), .IN8(~na473_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x45y95     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a475_4 ( .OUT(na475_2), .IN1(na135_1), .IN2(na448_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x44y99     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a476_1 ( .OUT(na476_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1136_1), .IN7(na25_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x48y94     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a477_1 ( .OUT(na477_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1), .IN8(na1526_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a477_2 ( .OUT(na477_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na477_1_i) );
// C_MX2b////      x48y91     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a478_1 ( .OUT(na478_1), .IN1(1'b1), .IN2(~na1441_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1173_1), .IN8(~na473_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x41y87     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a479_1 ( .OUT(na479_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na135_2), .IN6(na448_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y101     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a480_1 ( .OUT(na480_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na25_1), .IN8(na1138_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x49y94     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a481_1 ( .OUT(na481_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1), .IN8(na1527_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a481_2 ( .OUT(na481_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na481_1_i) );
// C_MX2b////      x49y91     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a482_1 ( .OUT(na482_1), .IN1(1'b1), .IN2(~na1441_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1174_1), .IN8(~na477_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y91     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a483_1 ( .OUT(na483_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na353_2), .IN6(~na448_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x45y101     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a484_1 ( .OUT(na484_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(1'b1), .IN7(na25_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x49y94     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a485_4 ( .OUT(na485_2_i), .IN1(na1528_1), .IN2(na470_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a485_5 ( .OUT(na485_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na485_2_i) );
// C_MX2b////      x47y91     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a486_1 ( .OUT(na486_1), .IN1(1'b1), .IN2(~na1441_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1175_1), .IN6(~na481_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x50y89     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a487_4 ( .OUT(na487_2), .IN1(~na1648_2), .IN2(na355_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x43y101     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a488_1 ( .OUT(na488_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na25_1), .IN8(na1143_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x49y93     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a489_4 ( .OUT(na489_2_i), .IN1(1'b1), .IN2(na470_2), .IN3(na1529_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a489_5 ( .OUT(na489_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na489_2_i) );
// C_MX2b////      x47y94     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a490_1 ( .OUT(na490_1), .IN1(1'b1), .IN2(~na1441_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1176_1), .IN6(~na485_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y89     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a491_1 ( .OUT(na491_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na448_2), .IN7(1'b1), .IN8(na309_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y90     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a492_1 ( .OUT(na492_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na448_2), .IN7(na497_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x41y99     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a493_4 ( .OUT(na493_2), .IN1(na1150_1), .IN2(1'b1), .IN3(na25_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x52y112     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a494_1 ( .OUT(na494_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1), .IN8(na1530_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a494_2 ( .OUT(na494_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na494_1_i) );
// C_MX2b////      x48y95     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a495_1 ( .OUT(na495_1), .IN1(1'b1), .IN2(na1441_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na379_2), .IN8(~na1177_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x48y89     80'h00_FE00_80_0000_0C08_FFC4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a497_4 ( .OUT(na497_2_i), .IN1(~na311_2), .IN2(na470_2), .IN3(1'b1), .IN4(na1532_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a497_5 ( .OUT(na497_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na497_2_i) );
// C_///AND*/D      x36y109     80'h00_FE00_80_0000_0C07_FF55
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a498_4 ( .OUT(na498_2_i), .IN1(~na1653_2), .IN2(1'b1), .IN3(~na844_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a498_5 ( .OUT(na498_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na498_2_i) );
// C_AND/D//AND/D      x21y116     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a499_1 ( .OUT(na499_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1178_1), .IN6(na663_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a499_2 ( .OUT(na499_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na499_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a499_4 ( .OUT(na499_2_i), .IN1(na1178_1), .IN2(na663_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a499_5 ( .OUT(na499_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na499_2_i) );
// C_AND/D//AND/D      x22y117     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a501_1 ( .OUT(na501_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na661_2), .IN6(na1178_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a501_2 ( .OUT(na501_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na501_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a501_4 ( .OUT(na501_2_i), .IN1(na661_1), .IN2(na1178_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a501_5 ( .OUT(na501_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na501_2_i) );
// C_AND/D//AND/D      x22y116     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a503_1 ( .OUT(na503_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1178_1), .IN6(na659_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a503_2 ( .OUT(na503_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na503_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a503_4 ( .OUT(na503_2_i), .IN1(na1178_1), .IN2(na659_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a503_5 ( .OUT(na503_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na503_2_i) );
// C_AND/D//AND/D      x24y116     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a505_1 ( .OUT(na505_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na656_2), .IN6(na1178_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a505_2 ( .OUT(na505_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na505_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a505_4 ( .OUT(na505_2_i), .IN1(na656_1), .IN2(na1178_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a505_5 ( .OUT(na505_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na505_2_i) );
// C_AND/D//AND/D      x23y114     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a507_1 ( .OUT(na507_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1178_1), .IN6(na654_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a507_2 ( .OUT(na507_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na507_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a507_4 ( .OUT(na507_2_i), .IN1(na1178_1), .IN2(na654_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a507_5 ( .OUT(na507_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na507_2_i) );
// C_AND/D//AND/D      x22y103     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a509_1 ( .OUT(na509_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1178_1), .IN6(na668_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a509_2 ( .OUT(na509_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na509_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a509_4 ( .OUT(na509_2_i), .IN1(na1178_1), .IN2(na668_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a509_5 ( .OUT(na509_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na509_2_i) );
// C_AND/D//AND/D      x22y108     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a511_1 ( .OUT(na511_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na670_2), .IN6(na1178_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a511_2 ( .OUT(na511_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na511_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a511_4 ( .OUT(na511_2_i), .IN1(na670_1), .IN2(na1178_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a511_5 ( .OUT(na511_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na511_2_i) );
// C_AND/D//AND/D      x24y105     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a513_1 ( .OUT(na513_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1178_1), .IN6(na672_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a513_2 ( .OUT(na513_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na513_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a513_4 ( .OUT(na513_2_i), .IN1(na1178_1), .IN2(na672_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a513_5 ( .OUT(na513_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na513_2_i) );
// C_AND/D//AND/D      x24y106     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a515_1 ( .OUT(na515_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na648_2), .IN6(na1178_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a515_2 ( .OUT(na515_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na515_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a515_4 ( .OUT(na515_2_i), .IN1(na648_1), .IN2(na1178_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a515_5 ( .OUT(na515_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na515_2_i) );
// C_AND/D//AND/D      x24y109     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a517_1 ( .OUT(na517_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1178_1), .IN6(na650_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a517_2 ( .OUT(na517_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na517_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a517_4 ( .OUT(na517_2_i), .IN1(na1178_1), .IN2(na650_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a517_5 ( .OUT(na517_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na517_2_i) );
// C_AND/D//AND/D      x23y111     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a519_1 ( .OUT(na519_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na652_2), .IN6(na1178_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a519_2 ( .OUT(na519_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na519_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a519_4 ( .OUT(na519_2_i), .IN1(na652_1), .IN2(na1178_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a519_5 ( .OUT(na519_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na519_2_i) );
// C_AND/D///      x23y101     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a522_1 ( .OUT(na522_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1178_1), .IN6(na657_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a522_2 ( .OUT(na522_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na522_1_i) );
// C_AND/D//AND/D      x24y104     80'h00_FE00_80_0000_0C88_F83A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a523_1 ( .OUT(na523_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1178_1), .IN6(na657_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a523_2 ( .OUT(na523_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na523_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a523_4 ( .OUT(na523_2_i), .IN1(na1178_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na523_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a523_5 ( .OUT(na523_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na523_2_i) );
// C_AND/D//AND/D      x24y103     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a525_1 ( .OUT(na525_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na666_2), .IN6(na1178_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a525_2 ( .OUT(na525_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na525_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a525_4 ( .OUT(na525_2_i), .IN1(na666_1), .IN2(na1178_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a525_5 ( .OUT(na525_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na525_2_i) );
// C_AND////      x44y101     80'h00_0018_00_0000_0888_3CC8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a526_1 ( .OUT(na526_1), .IN1(na1557_2), .IN2(na267_1), .IN3(1'b1), .IN4(na420_2), .IN5(1'b1), .IN6(na470_2), .IN7(1'b1),
                     .IN8(~na416_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x36y102     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a527_4 ( .OUT(na527_2), .IN1(na39_2), .IN2(na1559_2), .IN3(na250_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y98     80'h00_0018_00_0000_0888_AA4A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a528_1 ( .OUT(na528_1), .IN1(na23_1), .IN2(1'b1), .IN3(~na241_1), .IN4(na292_1), .IN5(na1363_2), .IN6(1'b1), .IN7(na44_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x32y111     80'h00_FE00_00_0000_0888_8C24
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a529_1 ( .OUT(na529_1_i), .IN1(~na1674_2), .IN2(na533_1), .IN3(na536_1), .IN4(~na1010_2), .IN5(1'b1), .IN6(na1654_2), .IN7(na536_2),
                     .IN8(na535_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a529_2 ( .OUT(na529_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na529_1_i) );
// C_AND////      x25y118     80'h00_0018_00_0000_0888_5111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a533_1 ( .OUT(na533_1), .IN1(~na1672_2), .IN2(~na1030_1), .IN3(~na1695_2), .IN4(~na741_1), .IN5(~na1673_2), .IN6(~na1026_2),
                     .IN7(~na747_1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x24y114     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a535_1 ( .OUT(na535_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1022_2), .IN6(~na1012_1), .IN7(~na1620_2),
                     .IN8(~na748_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a535_4 ( .OUT(na535_2), .IN1(~na1022_1), .IN2(~na1028_1), .IN3(~na743_1), .IN4(~na745_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x30y111     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a536_1 ( .OUT(na536_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1018_2), .IN6(~na1016_2), .IN7(~na759_1),
                     .IN8(~na761_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a536_4 ( .OUT(na536_2), .IN1(~na1018_1), .IN2(~na1016_1), .IN3(~na739_1), .IN4(~na757_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x38y112     80'h00_FE00_00_0000_0888_C844
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a537_1 ( .OUT(na537_1_i), .IN1(~na900_1), .IN2(na543_1), .IN3(~na847_1), .IN4(na544_1), .IN5(na541_1), .IN6(na543_2), .IN7(1'b1),
                     .IN8(na544_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a537_2 ( .OUT(na537_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na537_1_i) );
// C_AND////      x29y115     80'h00_0018_00_0000_0888_5111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a541_1 ( .OUT(na541_1), .IN1(~na1692_2), .IN2(~na920_1), .IN3(~na1694_2), .IN4(~na833_1), .IN5(~na1693_2), .IN6(~na916_1),
                     .IN7(~na839_1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x35y112     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a543_1 ( .OUT(na543_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na902_2), .IN6(~na912_2), .IN7(~na498_2), .IN8(~na840_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a543_4 ( .OUT(na543_2), .IN1(~na918_2), .IN2(~na912_1), .IN3(~na835_1), .IN4(~na837_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x38y110     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a544_1 ( .OUT(na544_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na906_2), .IN6(~na908_2), .IN7(~na851_1), .IN8(~na853_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a544_4 ( .OUT(na544_2), .IN1(~na906_1), .IN2(~na908_1), .IN3(~na831_1), .IN4(~na849_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x51y118     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a545_1 ( .OUT(na545_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na388_2), .IN7(na331_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x19y87     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a546_1 ( .OUT(na546_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na328_2), .IN6(na260_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x46y101     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a547_4 ( .OUT(na547_2), .IN1(na383_1), .IN2(1'b1), .IN3(na1032_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y96     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a548_1 ( .OUT(na548_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na383_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1033_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x46y100     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a549_4 ( .OUT(na549_2), .IN1(na383_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1034_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x45y96     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a550_1 ( .OUT(na550_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1035_1), .IN6(1'b1), .IN7(na1641_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x45y98     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a551_1 ( .OUT(na551_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na383_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1036_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x44y102     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a552_4 ( .OUT(na552_2), .IN1(na383_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1037_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x45y98     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a553_4 ( .OUT(na553_2), .IN1(na383_1), .IN2(na1039_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y100     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a554_4 ( .OUT(na554_2), .IN1(1'b1), .IN2(na922_1), .IN3(na250_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y99     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a555_4 ( .OUT(na555_2), .IN1(1'b1), .IN2(na1613_2), .IN3(na923_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y101     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a556_4 ( .OUT(na556_2), .IN1(1'b1), .IN2(1'b1), .IN3(na250_2), .IN4(na924_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x27y99     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a557_1 ( .OUT(na557_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na925_2), .IN7(na250_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x26y104     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a558_4 ( .OUT(na558_2), .IN1(1'b1), .IN2(na926_1), .IN3(na250_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x26y99     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a559_1 ( .OUT(na559_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na250_2), .IN8(na927_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x32y104     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a560_1 ( .OUT(na560_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na928_1), .IN6(1'b1), .IN7(na250_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x26y90     80'h00_0018_00_0040_0C09_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a576_1 ( .OUT(na576_1), .IN1(na1228_2), .IN2(1'b0), .IN3(1'b0), .IN4(na164_1), .IN5(na166_1), .IN6(1'b1), .IN7(~na167_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y93     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a577_1 ( .OUT(na577_1), .IN1(1'b1), .IN2(~na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1534_2), .IN8(na807_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D//OR/D      x39y94     80'h00_FE00_80_0000_0CEE_D05A
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a578_1 ( .OUT(na578_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na44_1), .IN8(na1535_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a578_2 ( .OUT(na578_1), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na578_1_i) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a578_4 ( .OUT(na578_2_i), .IN1(na1278_1), .IN2(1'b0), .IN3(~na44_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a578_5 ( .OUT(na578_2), .CLK(na1197_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na578_2_i) );
// C_MX4a////      x47y117     80'h00_0018_00_0040_0C09_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a579_1 ( .OUT(na579_1), .IN1(na1704_2), .IN2(1'b0), .IN3(1'b0), .IN4(na1138_1), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1143_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x45y109     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a580_1 ( .OUT(na580_1), .IN1(~na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1537_1), .IN8(na715_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D//OR/D      x45y102     80'h00_FE00_80_0000_0CEE_5CA3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a581_1 ( .OUT(na581_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1538_1), .IN7(~na1650_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a581_2 ( .OUT(na581_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na581_1_i) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a581_4 ( .OUT(na581_2_i), .IN1(1'b0), .IN2(~na470_2), .IN3(na1504_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a581_5 ( .OUT(na581_2), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na581_2_i) );
// C_ADDF2///ADDF2/      x33y98     80'h00_0078_00_0020_0C66_ACC5
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a582_1 ( .OUT(na582_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1116_2), .IN7(na241_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na583_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a582_4 ( .OUT(na582_2), .COUTY1(na582_4), .IN1(~na780_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1607_2), .IN5(1'b1), .IN6(na1116_2),
                     .IN7(na241_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na583_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x33y97     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a583_2 ( .OUT(na583_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a583_6 ( .COUTY1(na583_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na583_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x33y99     80'h00_0078_00_0020_0C66_C5A3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a604_1 ( .OUT(na604_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na780_2), .IN6(1'b1), .IN7(1'b1), .IN8(na270_2),
                     .CINX(1'b0), .CINY1(na582_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a604_4 ( .OUT(na604_2), .COUTY1(na604_4), .IN1(1'b1), .IN2(~na782_1), .IN3(na272_2), .IN4(1'b1), .IN5(~na780_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na270_2), .CINX(1'b0), .CINY1(na582_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x33y100     80'h00_0078_00_0020_0C66_C3C5
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a608_1 ( .OUT(na608_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na782_2), .IN7(1'b1), .IN8(na270_1),
                     .CINX(1'b0), .CINY1(na604_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a608_4 ( .OUT(na608_2), .COUTY1(na608_4), .IN1(~na785_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1608_2), .IN5(1'b1), .IN6(~na782_2),
                     .IN7(1'b1), .IN8(na270_1), .CINX(1'b0), .CINY1(na604_4), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x33y101     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a610_1 ( .OUT(na610_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0), .CINX(1'b0),
                     .CINY1(na608_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x39y103     80'h00_0078_00_0020_0C66_CA5A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a614_1 ( .OUT(na614_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na994_2), .IN6(1'b1), .IN7(1'b1), .IN8(na416_1),
                     .CINX(1'b0), .CINY1(na615_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a614_4 ( .OUT(na614_2), .COUTY1(na614_4), .IN1(na402_2), .IN2(1'b1), .IN3(~na691_1), .IN4(1'b1), .IN5(na994_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na416_1), .CINX(1'b0), .CINY1(na615_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x39y102     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a615_2 ( .OUT(na615_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a615_6 ( .COUTY1(na615_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na615_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x39y104     80'h00_0078_00_0020_0C66_5A3A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a636_1 ( .OUT(na636_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na412_2), .IN6(1'b1), .IN7(~na691_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na614_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a636_4 ( .OUT(na636_2), .COUTY1(na636_4), .IN1(na412_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na693_1), .IN5(na412_2), .IN6(1'b1),
                     .IN7(~na691_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na614_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x39y105     80'h00_0078_00_0020_0C66_3C5A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a640_1 ( .OUT(na640_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na410_1), .IN7(1'b1), .IN8(~na693_2),
                     .CINX(1'b0), .CINY1(na636_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a640_4 ( .OUT(na640_2), .COUTY1(na640_4), .IN1(na402_1), .IN2(1'b1), .IN3(~na696_1), .IN4(1'b1), .IN5(1'b1), .IN6(na410_1),
                     .IN7(1'b1), .IN8(~na693_2), .CINX(1'b0), .CINY1(na636_4), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x39y106     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a642_1 ( .OUT(na642_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0), .CINX(1'b0),
                     .CINY1(na640_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y107     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a648_1 ( .OUT(na648_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na515_2),
                     .CINX(1'b0), .CINY1(na672_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a648_4 ( .OUT(na648_2), .COUTY1(na648_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na515_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na515_2), .CINX(1'b0), .CINY1(na672_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y108     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a650_1 ( .OUT(na650_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na517_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na648_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a650_4 ( .OUT(na650_2), .COUTY1(na650_4), .IN1(1'b0), .IN2(1'b0), .IN3(na517_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na517_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na648_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y109     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a652_1 ( .OUT(na652_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na519_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na650_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a652_4 ( .OUT(na652_2), .COUTY1(na652_4), .IN1(na519_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na519_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na650_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y110     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a654_1 ( .OUT(na654_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na507_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na652_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a654_4 ( .OUT(na654_2), .COUTY1(na654_4), .IN1(1'b1), .IN2(na507_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na507_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na652_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y111     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a656_1 ( .OUT(na656_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na505_2),
                     .CINX(1'b0), .CINY1(na654_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a656_4 ( .OUT(na656_2), .COUTY1(na656_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na505_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na505_2), .CINX(1'b0), .CINY1(na654_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y102     80'h00_0078_00_0020_0C66_CAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a657_1 ( .OUT(na657_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na522_1), .IN6(1'b1), .IN7(1'b1), .IN8(na523_2),
                     .CINX(1'b0), .CINY1(na673_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a657_4 ( .OUT(na657_2), .COUTY1(na657_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na523_1), .IN5(na522_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na523_2), .CINX(1'b0), .CINY1(na673_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y112     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a659_1 ( .OUT(na659_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na503_2),
                     .CINX(1'b0), .CINY1(na656_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a659_4 ( .OUT(na659_2), .COUTY1(na659_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na503_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na503_2), .CINX(1'b0), .CINY1(na656_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y113     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a661_1 ( .OUT(na661_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na501_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na659_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a661_4 ( .OUT(na661_2), .COUTY1(na661_4), .IN1(1'b0), .IN2(1'b0), .IN3(na501_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na501_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na659_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y114     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a663_1 ( .OUT(na663_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na499_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na661_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a663_4 ( .OUT(na663_2), .IN1(1'b1), .IN2(na499_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na499_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na661_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y103     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a666_1 ( .OUT(na666_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na525_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na657_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a666_4 ( .OUT(na666_2), .COUTY1(na666_4), .IN1(1'b0), .IN2(1'b0), .IN3(na525_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na525_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na657_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y104     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a668_1 ( .OUT(na668_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na509_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na666_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a668_4 ( .OUT(na668_2), .COUTY1(na668_4), .IN1(1'b0), .IN2(1'b0), .IN3(na509_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na509_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na666_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y105     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a670_1 ( .OUT(na670_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na511_2),
                     .CINX(1'b0), .CINY1(na668_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a670_4 ( .OUT(na670_2), .COUTY1(na670_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na511_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na511_2), .CINX(1'b0), .CINY1(na668_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x21y106     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a672_1 ( .OUT(na672_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na513_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na670_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a672_4 ( .OUT(na672_2), .COUTY1(na672_4), .IN1(1'b0), .IN2(1'b0), .IN3(na513_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na513_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na670_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x21y101     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a673_2 ( .OUT(na673_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a673_6 ( .COUTY1(na673_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na673_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x41y101     80'h00_0078_00_0020_0C66_ACC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a675_1 ( .OUT(na675_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1639_2), .IN7(na331_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na684_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a675_4 ( .OUT(na675_2), .COUTY1(na675_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na367_1), .IN5(1'b1), .IN6(na1639_2),
                     .IN7(na331_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na684_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x41y102     80'h00_0078_00_0020_0C66_0AC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a677_1 ( .OUT(na677_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na372_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na675_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a677_4 ( .OUT(na677_2), .COUTY1(na677_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na177_2), .IN5(na372_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na675_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x41y103     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a679_1 ( .OUT(na679_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na182_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na677_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a679_4 ( .OUT(na679_2), .COUTY1(na679_4), .IN1(1'b0), .IN2(1'b0), .IN3(na179_2), .IN4(1'b1), .IN5(na182_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na677_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x41y104     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a681_1 ( .OUT(na681_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na184_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na679_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a681_4 ( .OUT(na681_2), .COUTY1(na681_4), .IN1(1'b0), .IN2(1'b0), .IN3(na17_2), .IN4(1'b1), .IN5(1'b1), .IN6(na184_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na679_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x41y105     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a683_1 ( .OUT(na683_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na11_2),
                     .CINX(1'b0), .CINY1(na681_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a683_4 ( .OUT(na683_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na19_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na11_2),
                     .CINX(1'b0), .CINY1(na681_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x41y100     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a684_2 ( .OUT(na684_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a684_6 ( .COUTY1(na684_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na684_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x37y99     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a685_1 ( .OUT(na685_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na402_2), .IN6(1'b1), .IN7(1'b1), .IN8(na416_1),
                     .CINX(1'b0), .CINY1(na690_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a685_4 ( .OUT(na685_2), .COUTY1(na685_4), .IN1(na412_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na402_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na416_1), .CINX(1'b0), .CINY1(na690_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x37y100     80'h00_0078_00_0020_0C66_0A0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a687_1 ( .OUT(na687_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na412_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na685_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a687_4 ( .OUT(na687_2), .COUTY1(na687_4), .IN1(1'b1), .IN2(na410_1), .IN3(1'b0), .IN4(1'b0), .IN5(na412_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na685_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x37y101     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a689_1 ( .OUT(na689_1), .IN1(na402_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na687_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x37y98     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a690_2 ( .OUT(na690_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a690_6 ( .COUTY1(na690_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na690_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x38y105     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a691_1 ( .OUT(na691_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na994_2), .IN6(1'b1), .IN7(1'b1), .IN8(na993_1),
                     .CINX(1'b0), .CINY1(na695_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a691_4 ( .OUT(na691_2), .COUTY1(na691_4), .IN1(na994_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na994_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na993_1), .CINX(1'b0), .CINY1(na695_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y106     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a693_1 ( .OUT(na693_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na996_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na691_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a693_4 ( .OUT(na693_2), .COUTY1(na693_4), .IN1(na996_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na996_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na691_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x38y104     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a695_2 ( .OUT(na695_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a695_6 ( .COUTY1(na695_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na695_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x38y107     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a696_1 ( .OUT(na696_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0), .CINX(1'b0),
                     .CINY1(na693_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y90     80'h00_0078_00_0020_0C66_CA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a697_1 ( .OUT(na697_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na353_2), .IN6(1'b1), .IN7(1'b1), .IN8(na309_2),
                     .CINX(1'b0), .CINY1(na702_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a697_4 ( .OUT(na697_2), .COUTY1(na697_4), .IN1(1'b1), .IN2(na355_2), .IN3(1'b0), .IN4(1'b0), .IN5(na353_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na309_2), .CINX(1'b0), .CINY1(na702_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y91     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a699_1 ( .OUT(na699_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na353_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na697_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a699_4 ( .OUT(na699_2), .COUTY1(na699_4), .IN1(1'b0), .IN2(1'b0), .IN3(na324_2), .IN4(1'b1), .IN5(na353_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na697_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x51y92     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a701_1 ( .OUT(na701_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na309_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na699_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x51y89     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a702_2 ( .OUT(na702_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a702_6 ( .COUTY1(na702_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na702_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x45y87     80'h00_0078_00_0020_0C66_CC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a703_1 ( .OUT(na703_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1635_2), .IN7(1'b1), .IN8(na343_1),
                     .CINX(1'b0), .CINY1(na709_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a703_4 ( .OUT(na703_2), .COUTY1(na703_4), .IN1(1'b1), .IN2(na337_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1635_2),
                     .IN7(1'b1), .IN8(na343_1), .CINX(1'b0), .CINY1(na709_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x45y88     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a705_1 ( .OUT(na705_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na497_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na703_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a705_4 ( .OUT(na705_2), .COUTY1(na705_4), .IN1(1'b1), .IN2(na337_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na497_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na703_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x45y89     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a707_1 ( .OUT(na707_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na135_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na705_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a707_4 ( .OUT(na707_2), .IN1(na135_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na135_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na705_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x45y86     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a709_2 ( .OUT(na709_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a709_6 ( .COUTY1(na709_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na709_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x48y104     80'h00_0078_00_0020_0C66_FAFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a711_1 ( .OUT(na711_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na459_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na736_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a711_4 ( .OUT(na711_2), .COUTY1(na711_4), .IN1(na456_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na459_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na736_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y105     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a713_1 ( .OUT(na713_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na453_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na711_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a713_4 ( .OUT(na713_2), .COUTY1(na713_4), .IN1(1'b1), .IN2(na287_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na453_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na711_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y106     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a715_1 ( .OUT(na715_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na581_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na713_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a715_4 ( .OUT(na715_2), .COUTY1(na715_4), .IN1(1'b1), .IN2(na581_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na581_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na713_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y107     80'h00_0078_00_0020_0C66_FCAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a717_1 ( .OUT(na717_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na441_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na715_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a717_4 ( .OUT(na717_2), .COUTY1(na717_4), .IN1(1'b1), .IN2(1'b1), .IN3(na282_2), .IN4(1'b1), .IN5(1'b1), .IN6(na441_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na715_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y108     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a719_1 ( .OUT(na719_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na436_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na717_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a719_4 ( .OUT(na719_2), .COUTY1(na719_4), .IN1(1'b1), .IN2(na436_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na436_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na717_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y99     80'h00_0078_00_0020_0C66_CAFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a720_1 ( .OUT(na720_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na391_2), .IN6(1'b1), .IN7(1'b1), .IN8(na418_2),
                     .CINX(1'b0), .CINY1(na737_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a720_4 ( .OUT(na720_2), .COUTY1(na720_4), .IN1(na391_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na391_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na418_2), .CINX(1'b0), .CINY1(na737_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y109     80'h00_0078_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a722_1 ( .OUT(na722_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na432_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na719_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a722_4 ( .OUT(na722_2), .COUTY1(na722_4), .IN1(1'b1), .IN2(1'b1), .IN3(na432_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na432_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na719_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y110     80'h00_0078_00_0020_0C66_CFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a724_1 ( .OUT(na724_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na427_2),
                     .CINX(1'b0), .CINY1(na722_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a724_4 ( .OUT(na724_2), .COUTY1(na724_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na427_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na427_2), .CINX(1'b0), .CINY1(na722_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y111     80'h00_0078_00_0020_0C66_CFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a726_1 ( .OUT(na726_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na421_2),
                     .CINX(1'b0), .CINY1(na724_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a726_4 ( .OUT(na726_2), .COUTY1(na726_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na421_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na421_2), .CINX(1'b0), .CINY1(na724_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x48y112     80'h00_0018_00_0010_0666_00FA
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a728_1 ( .OUT(na728_1), .IN1(na265_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na726_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y100     80'h00_0078_00_0020_0C66_FACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a730_1 ( .OUT(na730_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na385_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na720_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a730_4 ( .OUT(na730_2), .COUTY1(na730_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na111_2), .IN5(na385_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na720_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y101     80'h00_0078_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a732_1 ( .OUT(na732_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na80_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na730_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a732_4 ( .OUT(na732_2), .COUTY1(na732_4), .IN1(1'b1), .IN2(1'b1), .IN3(na80_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na80_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na730_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y102     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a734_1 ( .OUT(na734_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na66_1),
                     .CINX(1'b0), .CINY1(na732_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a734_4 ( .OUT(na734_2), .COUTY1(na734_4), .IN1(na465_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na66_1), .CINX(1'b0), .CINY1(na732_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y103     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a736_1 ( .OUT(na736_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na461_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na734_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a736_4 ( .OUT(na736_2), .COUTY1(na736_4), .IN1(1'b1), .IN2(na461_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na461_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na734_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x48y98     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a737_2 ( .OUT(na737_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a737_6 ( .COUTY1(na737_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na737_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x26y111     80'h00_F660_00_0020_0C66_AFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a739_1 ( .OUT(na739_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na739_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na761_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a739_2 ( .OUT(na739_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na739_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a739_4 ( .OUT(na739_2), .COUTY1(na739_4), .IN1(na1018_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na739_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na761_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x26y112     80'h00_F660_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a741_1 ( .OUT(na741_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na741_1),
                     .CINX(1'b0), .CINY1(na739_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a741_2 ( .OUT(na741_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na741_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a741_4 ( .OUT(na741_2), .COUTY1(na741_4), .IN1(na1022_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na741_1), .CINX(1'b0), .CINY1(na739_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x26y113     80'h00_F660_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a743_1 ( .OUT(na743_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na743_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na741_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a743_2 ( .OUT(na743_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na743_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a743_4 ( .OUT(na743_2), .COUTY1(na743_4), .IN1(1'b1), .IN2(na1030_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na743_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na741_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x26y114     80'h00_F660_00_0020_0C66_CFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a745_1 ( .OUT(na745_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na745_1),
                     .CINX(1'b0), .CINY1(na743_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a745_2 ( .OUT(na745_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na745_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a745_4 ( .OUT(na745_2), .COUTY1(na745_4), .IN1(1'b1), .IN2(na1026_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na745_1), .CINX(1'b0), .CINY1(na743_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x26y115     80'h00_F660_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a747_1 ( .OUT(na747_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na747_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na745_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a747_2 ( .OUT(na747_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na747_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a747_4 ( .OUT(na747_2), .COUTY1(na747_4), .IN1(1'b1), .IN2(na1028_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na747_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na745_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x26y106     80'h00_F660_00_0020_0C66_CACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a748_1 ( .OUT(na748_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1022_2), .IN6(1'b1), .IN7(1'b1), .IN8(na748_1),
                     .CINX(1'b0), .CINY1(na762_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a748_2 ( .OUT(na748_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na748_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a748_4 ( .OUT(na748_2), .COUTY1(na748_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1010_2), .IN5(na1022_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na748_1), .CINX(1'b0), .CINY1(na762_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x26y116     80'h00_F660_00_0020_0C66_CFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a750_1 ( .OUT(na750_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na750_1),
                     .CINX(1'b0), .CINY1(na747_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a750_2 ( .OUT(na750_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na750_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a750_4 ( .OUT(na750_2), .COUTY1(na750_4), .IN1(1'b1), .IN2(na1030_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na750_1), .CINX(1'b0), .CINY1(na747_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x26y117     80'h00_F660_00_0020_0C66_AFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a752_1 ( .OUT(na752_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na752_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na750_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a752_2 ( .OUT(na752_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na752_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a752_4 ( .OUT(na752_2), .IN1(na291_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na752_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na750_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x26y107     80'h00_F660_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a755_1 ( .OUT(na755_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na755_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na748_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a755_2 ( .OUT(na755_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na755_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a755_4 ( .OUT(na755_2), .COUTY1(na755_4), .IN1(1'b1), .IN2(na1012_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na755_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na748_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x26y108     80'h00_F660_00_0020_0C66_CFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a757_1 ( .OUT(na757_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na757_1),
                     .CINX(1'b0), .CINY1(na755_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a757_2 ( .OUT(na757_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na757_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a757_4 ( .OUT(na757_2), .COUTY1(na757_4), .IN1(1'b1), .IN2(na1016_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na757_1), .CINX(1'b0), .CINY1(na755_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x26y109     80'h00_F660_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a759_1 ( .OUT(na759_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na759_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na757_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a759_2 ( .OUT(na759_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na759_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a759_4 ( .OUT(na759_2), .COUTY1(na759_4), .IN1(1'b1), .IN2(na1016_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na759_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na757_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x26y110     80'h00_F660_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a761_1 ( .OUT(na761_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na761_1),
                     .CINX(1'b0), .CINY1(na759_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a761_2 ( .OUT(na761_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na761_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a761_4 ( .OUT(na761_2), .COUTY1(na761_4), .IN1(na1018_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na761_1), .CINX(1'b0), .CINY1(na759_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x26y105     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a762_2 ( .OUT(na762_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a762_6 ( .COUTY1(na762_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na762_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x22y91     80'h00_0078_00_0020_0C66_CAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a764_1 ( .OUT(na764_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na328_2), .IN6(1'b1), .IN7(1'b1), .IN8(na323_2),
                     .CINX(1'b0), .CINY1(na773_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a764_4 ( .OUT(na764_2), .COUTY1(na764_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na323_1), .IN5(na328_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na323_2), .CINX(1'b0), .CINY1(na773_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x22y92     80'h00_0078_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a766_1 ( .OUT(na766_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na322_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na764_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a766_4 ( .OUT(na766_2), .COUTY1(na766_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na139_2), .IN5(1'b0), .IN6(1'b0), .IN7(na322_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na764_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x22y93     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a768_1 ( .OUT(na768_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na137_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na766_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a768_4 ( .OUT(na768_2), .COUTY1(na768_4), .IN1(1'b0), .IN2(1'b0), .IN3(na141_2), .IN4(1'b1), .IN5(na137_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na766_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x22y94     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a770_1 ( .OUT(na770_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na377_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na768_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a770_4 ( .OUT(na770_2), .COUTY1(na770_4), .IN1(1'b0), .IN2(1'b0), .IN3(na375_2), .IN4(1'b1), .IN5(1'b1), .IN6(na377_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na768_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x22y95     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a772_1 ( .OUT(na772_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na155_2),
                     .CINX(1'b0), .CINY1(na770_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a772_4 ( .OUT(na772_2), .IN1(na258_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na155_2),
                     .CINX(1'b0), .CINY1(na770_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x22y90     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a773_2 ( .OUT(na773_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a773_6 ( .COUTY1(na773_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na773_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x33y107     80'h00_0078_00_0020_0C66_ACC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a774_1 ( .OUT(na774_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na219_1), .IN7(na241_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na779_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a774_4 ( .OUT(na774_2), .COUTY1(na774_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na270_2), .IN5(1'b1), .IN6(na219_1), .IN7(na241_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na779_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x33y108     80'h00_0078_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a776_1 ( .OUT(na776_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na272_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na774_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a776_4 ( .OUT(na776_2), .COUTY1(na776_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na270_1), .IN5(1'b0), .IN6(1'b0), .IN7(na272_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na774_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x33y109     80'h00_0018_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a778_1 ( .OUT(na778_1), .IN1(1'b1), .IN2(na219_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na776_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x33y106     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a779_2 ( .OUT(na779_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a779_6 ( .COUTY1(na779_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na779_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x35y99     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a780_1 ( .OUT(na780_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1116_2), .IN7(na1115_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na784_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a780_4 ( .OUT(na780_2), .COUTY1(na780_4), .IN1(1'b1), .IN2(na1116_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1116_2),
                     .IN7(na1115_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na784_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x35y100     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a782_1 ( .OUT(na782_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1118_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na780_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a782_4 ( .OUT(na782_2), .COUTY1(na782_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1118_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1118_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na780_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x35y98     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a784_2 ( .OUT(na784_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a784_6 ( .COUTY1(na784_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na784_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x35y101     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a785_1 ( .OUT(na785_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0), .CINX(1'b0),
                     .CINY1(na782_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x22y110     80'h00_0078_00_0020_0C66_AAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a786_1 ( .OUT(na786_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na231_1), .IN6(1'b1), .IN7(na314_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na793_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a786_4 ( .OUT(na786_2), .COUTY1(na786_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na318_1), .IN5(na231_1), .IN6(1'b1), .IN7(na314_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na793_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x22y111     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a788_1 ( .OUT(na788_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na316_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na786_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a788_4 ( .OUT(na788_2), .COUTY1(na788_4), .IN1(1'b0), .IN2(1'b0), .IN3(na314_1), .IN4(1'b1), .IN5(1'b1), .IN6(na316_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na786_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x22y112     80'h00_0078_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a790_1 ( .OUT(na790_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na316_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na788_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a790_4 ( .OUT(na790_2), .COUTY1(na790_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na318_2), .IN5(1'b1), .IN6(na316_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na788_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x22y113     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a792_1 ( .OUT(na792_1), .IN1(na231_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na790_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x22y109     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a793_2 ( .OUT(na793_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a793_6 ( .COUTY1(na793_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na793_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x28y110     80'h00_0078_00_0020_0C66_CAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a794_1 ( .OUT(na794_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na299_2), .IN6(1'b1), .IN7(1'b1), .IN8(na300_2),
                     .CINX(1'b0), .CINY1(na801_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a794_4 ( .OUT(na794_2), .COUTY1(na794_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na300_1), .IN5(na299_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na300_2), .CINX(1'b0), .CINY1(na801_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x28y111     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a796_1 ( .OUT(na796_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na299_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na794_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a796_4 ( .OUT(na796_2), .COUTY1(na796_4), .IN1(na297_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na299_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na794_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x28y112     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a798_1 ( .OUT(na798_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na298_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na796_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a798_4 ( .OUT(na798_2), .COUTY1(na798_4), .IN1(na297_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na298_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na796_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x28y113     80'h00_0018_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a800_1 ( .OUT(na800_1), .IN1(1'b1), .IN2(na293_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na798_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x28y109     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a801_2 ( .OUT(na801_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a801_6 ( .COUTY1(na801_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na801_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x36y92     80'h00_0078_00_0020_0C66_FAFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a803_1 ( .OUT(na803_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na92_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na828_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a803_4 ( .OUT(na803_2), .COUTY1(na803_4), .IN1(1'b1), .IN2(na95_1), .IN3(1'b1), .IN4(1'b1), .IN5(na92_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na828_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y93     80'h00_0078_00_0020_0C66_FACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a805_1 ( .OUT(na805_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na99_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na803_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a805_4 ( .OUT(na805_2), .COUTY1(na805_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na102_1), .IN5(na99_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na803_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y94     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a807_1 ( .OUT(na807_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na578_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na805_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a807_4 ( .OUT(na807_2), .COUTY1(na807_4), .IN1(1'b1), .IN2(na578_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na578_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na805_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y95     80'h00_0078_00_0020_0C66_FCCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a809_1 ( .OUT(na809_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na117_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na807_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a809_4 ( .OUT(na809_2), .COUTY1(na809_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na121_2), .IN5(1'b1), .IN6(na117_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na807_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y96     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a811_1 ( .OUT(na811_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na51_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na809_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a811_4 ( .OUT(na811_2), .COUTY1(na811_4), .IN1(1'b1), .IN2(na51_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na51_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na809_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y87     80'h00_0078_00_0020_0C66_CCCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a812_1 ( .OUT(na812_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na229_2), .IN7(1'b1), .IN8(na131_2),
                     .CINX(1'b0), .CINY1(na829_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a812_4 ( .OUT(na812_2), .COUTY1(na812_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na131_1), .IN5(1'b1), .IN6(na229_2), .IN7(1'b1),
                     .IN8(na131_2), .CINX(1'b0), .CINY1(na829_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y97     80'h00_0078_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a814_1 ( .OUT(na814_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na63_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na811_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a814_4 ( .OUT(na814_2), .COUTY1(na814_4), .IN1(1'b1), .IN2(1'b1), .IN3(na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na63_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na811_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y98     80'h00_0078_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a816_1 ( .OUT(na816_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na263_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na814_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a816_4 ( .OUT(na816_2), .COUTY1(na816_4), .IN1(1'b1), .IN2(1'b1), .IN3(na263_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na263_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na814_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y99     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a818_1 ( .OUT(na818_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na227_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na816_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a818_4 ( .OUT(na818_2), .COUTY1(na818_4), .IN1(1'b1), .IN2(na227_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na227_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na816_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x36y100     80'h00_0018_00_0010_0666_00FC
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a820_1 ( .OUT(na820_1), .IN1(1'b1), .IN2(na256_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na818_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y88     80'h00_0078_00_0020_0C66_FCAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a822_1 ( .OUT(na822_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na133_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na812_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a822_4 ( .OUT(na822_2), .COUTY1(na822_4), .IN1(1'b1), .IN2(1'b1), .IN3(na74_2), .IN4(1'b1), .IN5(1'b1), .IN6(na133_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na812_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y89     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a824_1 ( .OUT(na824_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na78_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na822_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a824_4 ( .OUT(na824_2), .COUTY1(na824_4), .IN1(1'b1), .IN2(na78_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na78_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na822_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y90     80'h00_0078_00_0020_0C66_FACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a826_1 ( .OUT(na826_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na224_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na824_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a826_4 ( .OUT(na826_2), .COUTY1(na826_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na83_2), .IN5(na224_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na824_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y91     80'h00_0078_00_0020_0C66_CFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a828_1 ( .OUT(na828_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na89_2),
                     .CINX(1'b0), .CINY1(na826_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a828_4 ( .OUT(na828_2), .COUTY1(na828_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na89_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na89_2), .CINX(1'b0), .CINY1(na826_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x36y86     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a829_2 ( .OUT(na829_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a829_6 ( .COUTY1(na829_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na829_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x34y109     80'h00_F660_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a831_1 ( .OUT(na831_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na831_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na853_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a831_2 ( .OUT(na831_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na831_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a831_4 ( .OUT(na831_2), .COUTY1(na831_4), .IN1(1'b1), .IN2(na908_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na831_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na853_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y110     80'h00_F660_00_0020_0C66_CFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a833_1 ( .OUT(na833_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na833_1),
                     .CINX(1'b0), .CINY1(na831_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a833_2 ( .OUT(na833_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na833_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a833_4 ( .OUT(na833_2), .COUTY1(na833_4), .IN1(1'b1), .IN2(na912_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na833_1), .CINX(1'b0), .CINY1(na831_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y111     80'h00_F660_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a835_1 ( .OUT(na835_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na835_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na833_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a835_2 ( .OUT(na835_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na835_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a835_4 ( .OUT(na835_2), .COUTY1(na835_4), .IN1(1'b1), .IN2(na920_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na835_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na833_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y112     80'h00_F660_00_0020_0C66_CFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a837_1 ( .OUT(na837_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na837_1),
                     .CINX(1'b0), .CINY1(na835_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a837_2 ( .OUT(na837_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na837_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a837_4 ( .OUT(na837_2), .COUTY1(na837_4), .IN1(1'b1), .IN2(na916_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na837_1), .CINX(1'b0), .CINY1(na835_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y113     80'h00_F660_00_0020_0C66_AFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a839_1 ( .OUT(na839_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na839_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na837_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a839_2 ( .OUT(na839_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na839_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a839_4 ( .OUT(na839_2), .COUTY1(na839_4), .IN1(na918_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na839_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na837_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y104     80'h00_F660_00_0020_0C66_CCFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a840_1 ( .OUT(na840_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na912_2), .IN7(1'b1), .IN8(na840_1),
                     .CINX(1'b0), .CINY1(na1207_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a840_2 ( .OUT(na840_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na840_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a840_4 ( .OUT(na840_2), .COUTY1(na840_4), .IN1(na900_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na912_2), .IN7(1'b1),
                     .IN8(na840_1), .CINX(1'b0), .CINY1(na1207_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y114     80'h00_F660_00_0020_0C66_CFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a842_1 ( .OUT(na842_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na842_1),
                     .CINX(1'b0), .CINY1(na839_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a842_2 ( .OUT(na842_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na842_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a842_4 ( .OUT(na842_2), .COUTY1(na842_4), .IN1(1'b1), .IN2(na920_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na842_1), .CINX(1'b0), .CINY1(na839_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y115     80'h00_F660_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a844_1 ( .OUT(na844_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na844_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na842_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a844_2 ( .OUT(na844_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na844_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a844_4 ( .OUT(na844_2), .IN1(1'b1), .IN2(1'b1), .IN3(na498_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na844_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na842_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y105     80'h00_F660_00_0020_0C66_AFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a847_1 ( .OUT(na847_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na847_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na840_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a847_2 ( .OUT(na847_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na847_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a847_4 ( .OUT(na847_2), .COUTY1(na847_4), .IN1(na902_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na847_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na840_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y106     80'h00_F660_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a849_1 ( .OUT(na849_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na849_1),
                     .CINX(1'b0), .CINY1(na847_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a849_2 ( .OUT(na849_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na849_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a849_4 ( .OUT(na849_2), .COUTY1(na849_4), .IN1(na906_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na849_1), .CINX(1'b0), .CINY1(na847_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y107     80'h00_F660_00_0020_0C66_AFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a851_1 ( .OUT(na851_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na851_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na849_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a851_2 ( .OUT(na851_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na851_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a851_4 ( .OUT(na851_2), .COUTY1(na851_4), .IN1(na906_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na851_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na849_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y108     80'h00_F660_00_0020_0C66_CFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a853_1 ( .OUT(na853_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na853_1),
                     .CINX(1'b0), .CINY1(na851_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a853_2 ( .OUT(na853_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na853_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a853_4 ( .OUT(na853_2), .COUTY1(na853_4), .IN1(1'b1), .IN2(na908_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na853_1), .CINX(1'b0), .CINY1(na851_4), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x35y109     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a900_1 ( .OUT(na900_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na840_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a900_2 ( .OUT(na900_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na900_1_i) );
// C_///AND/D      x37y109     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a902_4 ( .OUT(na902_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na847_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a902_5 ( .OUT(na902_2), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na902_2_i) );
// C_AND/D//AND/D      x37y111     80'h00_F600_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a906_1 ( .OUT(na906_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na851_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a906_2 ( .OUT(na906_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na906_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a906_4 ( .OUT(na906_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na849_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a906_5 ( .OUT(na906_2), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na906_2_i) );
// C_AND/D//AND/D      x37y112     80'h00_F600_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a908_1 ( .OUT(na908_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na853_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a908_2 ( .OUT(na908_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na908_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a908_4 ( .OUT(na908_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na831_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a908_5 ( .OUT(na908_2), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na908_2_i) );
// C_AND/D//AND/D      x39y110     80'h00_F600_80_0000_0C88_CFF3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a912_1 ( .OUT(na912_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na833_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a912_2 ( .OUT(na912_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na912_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a912_4 ( .OUT(na912_2_i), .IN1(1'b1), .IN2(~na912_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a912_5 ( .OUT(na912_2), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na912_2_i) );
// C_AND/D///      x29y114     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a916_1 ( .OUT(na916_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na837_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a916_2 ( .OUT(na916_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na916_1_i) );
// C_///AND/D      x27y115     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a918_4 ( .OUT(na918_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na839_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a918_5 ( .OUT(na918_2), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na918_2_i) );
// C_AND/D//AND/D      x29y116     80'h00_F600_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a920_1 ( .OUT(na920_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na842_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a920_2 ( .OUT(na920_1), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na920_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a920_4 ( .OUT(na920_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na835_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a920_5 ( .OUT(na920_2), .CLK(na1197_2), .EN(~na498_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na920_2_i) );
// C_AND/D///      x31y100     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a922_1 ( .OUT(na922_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na167_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a922_2 ( .OUT(na922_1), .CLK(na1197_2), .EN(na528_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na922_1_i) );
// C_///AND/D      x30y99     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a923_4 ( .OUT(na923_2_i), .IN1(1'b1), .IN2(na160_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a923_5 ( .OUT(na923_2), .CLK(na1197_2), .EN(na528_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na923_2_i) );
// C_///AND/D      x30y100     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a924_4 ( .OUT(na924_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na164_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a924_5 ( .OUT(na924_2), .CLK(na1197_2), .EN(na528_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na924_2_i) );
// C_///AND/D      x29y98     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a925_4 ( .OUT(na925_2_i), .IN1(na166_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a925_5 ( .OUT(na925_2), .CLK(na1197_2), .EN(na528_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na925_2_i) );
// C_AND/D///      x29y98     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a926_1 ( .OUT(na926_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na167_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a926_2 ( .OUT(na926_1), .CLK(na1197_2), .EN(na528_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na926_1_i) );
// C_///AND/D      x24y98     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a927_4 ( .OUT(na927_2_i), .IN1(na170_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a927_5 ( .OUT(na927_2), .CLK(na1197_2), .EN(na528_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na927_2_i) );
// C_AND/D///      x27y101     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a928_1 ( .OUT(na928_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na171_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a928_2 ( .OUT(na928_1), .CLK(na1197_2), .EN(na528_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na928_1_i) );
// C_///AND/D      x22y102     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a929_4 ( .OUT(na929_2_i), .IN1(1'b1), .IN2(na173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a929_5 ( .OUT(na929_2), .CLK(na1197_2), .EN(na528_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na929_2_i) );
// C_AND/D///      x42y110     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a993_1 ( .OUT(na993_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1136_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a993_2 ( .OUT(na993_1), .CLK(na1197_1), .EN(na400_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na993_1_i) );
// C_AND/D//AND/D      x41y109     80'h00_FA00_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a994_1 ( .OUT(na994_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1138_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a994_2 ( .OUT(na994_1), .CLK(na1197_1), .EN(na400_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na994_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a994_4 ( .OUT(na994_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1133_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a994_5 ( .OUT(na994_2), .CLK(na1197_1), .EN(na400_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na994_2_i) );
// C_AND/D//AND/D      x41y111     80'h00_FA00_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a996_1 ( .OUT(na996_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a996_2 ( .OUT(na996_1), .CLK(na1197_1), .EN(na400_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na996_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a996_4 ( .OUT(na996_2_i), .IN1(na1141_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a996_5 ( .OUT(na996_2), .CLK(na1197_1), .EN(na400_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na996_2_i) );
// C_///AND/D      x30y108     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1010_4 ( .OUT(na1010_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na748_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1010_5 ( .OUT(na1010_2), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1010_2_i) );
// C_AND/D///      x27y110     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1012_1 ( .OUT(na1012_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na755_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1012_2 ( .OUT(na1012_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1012_1_i) );
// C_AND/D//AND/D      x27y112     80'h00_F600_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1016_1 ( .OUT(na1016_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na759_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1016_2 ( .OUT(na1016_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1016_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1016_4 ( .OUT(na1016_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na757_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1016_5 ( .OUT(na1016_2), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1016_2_i) );
// C_AND/D//AND/D      x23y113     80'h00_F600_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1018_1 ( .OUT(na1018_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na761_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a1018_2 ( .OUT(na1018_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1018_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1018_4 ( .OUT(na1018_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na739_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a1018_5 ( .OUT(na1018_2), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1018_2_i) );
// C_AND/D//AND/D      x23y115     80'h00_F600_80_0000_0C88_CFF5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1022_1 ( .OUT(na1022_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na741_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1022_2 ( .OUT(na1022_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1022_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1022_4 ( .OUT(na1022_2_i), .IN1(~na1022_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1022_5 ( .OUT(na1022_2), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1022_2_i) );
// C_///AND/D      x27y118     80'h00_F600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1026_4 ( .OUT(na1026_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na745_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a1026_5 ( .OUT(na1026_2), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1026_2_i) );
// C_AND/D///      x21y118     80'h00_F600_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1028_1 ( .OUT(na1028_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na747_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a1028_2 ( .OUT(na1028_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1028_1_i) );
// C_AND/D//AND/D      x23y118     80'h00_F600_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1030_1 ( .OUT(na1030_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na750_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1030_2 ( .OUT(na1030_1), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1030_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1030_4 ( .OUT(na1030_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na743_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1030_5 ( .OUT(na1030_2), .CLK(na1197_1), .EN(~na291_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1030_2_i) );
// C_///AND/D      x42y117     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1032_4 ( .OUT(na1032_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1133_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1032_5 ( .OUT(na1032_2), .CLK(na1197_1), .EN(na526_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1032_2_i) );
// C_AND/D///      x44y108     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1033_1 ( .OUT(na1033_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1136_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1033_2 ( .OUT(na1033_1), .CLK(na1197_1), .EN(na526_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1033_1_i) );
// C_///AND/D      x44y112     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1034_4 ( .OUT(na1034_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1138_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1034_5 ( .OUT(na1034_2), .CLK(na1197_1), .EN(na526_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1034_2_i) );
// C_AND/D///      x43y107     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1035_1 ( .OUT(na1035_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1035_2 ( .OUT(na1035_1), .CLK(na1197_1), .EN(na526_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1035_1_i) );
// C_AND/D///      x46y108     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1036_1 ( .OUT(na1036_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1036_2 ( .OUT(na1036_1), .CLK(na1197_1), .EN(na526_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1036_1_i) );
// C_AND/D///      x42y106     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1037_1 ( .OUT(na1037_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1146_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1037_2 ( .OUT(na1037_1), .CLK(na1197_1), .EN(na526_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1037_1_i) );
// C_///AND/D      x41y98     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1038_4 ( .OUT(na1038_2_i), .IN1(na1147_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1038_5 ( .OUT(na1038_2), .CLK(na1197_1), .EN(na526_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1038_2_i) );
// C_AND/D///      x39y100     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1039_1 ( .OUT(na1039_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1150_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1039_2 ( .OUT(na1039_1), .CLK(na1197_1), .EN(na526_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1039_1_i) );
// C_///AND/D      x42y97     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1115_4 ( .OUT(na1115_2_i), .IN1(1'b1), .IN2(na160_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1115_5 ( .OUT(na1115_2), .CLK(na1197_2), .EN(na527_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1115_2_i) );
// C_AND/D//AND/D      x33y104     80'h00_FA00_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1116_1 ( .OUT(na1116_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na164_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1116_2 ( .OUT(na1116_1), .CLK(na1197_2), .EN(na527_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1116_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1116_4 ( .OUT(na1116_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na167_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1116_5 ( .OUT(na1116_2), .CLK(na1197_2), .EN(na527_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1116_2_i) );
// C_AND/D//AND/D      x32y101     80'h00_FA00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1118_1 ( .OUT(na1118_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na167_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1118_2 ( .OUT(na1118_1), .CLK(na1197_2), .EN(na527_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1118_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1118_4 ( .OUT(na1118_2_i), .IN1(na166_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1118_5 ( .OUT(na1118_2), .CLK(na1197_2), .EN(na527_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1118_2_i) );
// C_MX4b////      x33y112     80'h00_0018_00_0040_0A50_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1122_1 ( .OUT(na1122_1), .IN1(~na8_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1_2), .IN5(na778_1), .IN6(1'b0), .IN7(na1681_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x32y93     80'h00_0018_00_0040_0AF8_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1123_1 ( .OUT(na1123_1), .IN1(1'b1), .IN2(na377_1), .IN3(na375_1), .IN4(1'b1), .IN5(na152_1), .IN6(na153_1), .IN7(na154_1),
                      .IN8(~na151_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x24y90     80'h00_0018_00_0040_0AF0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1124_1 ( .OUT(na1124_1), .IN1(1'b1), .IN2(~na377_1), .IN3(~na375_1), .IN4(1'b1), .IN5(na159_1), .IN6(na143_1), .IN7(na158_2),
                      .IN8(na148_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x29y88     80'h00_0018_00_0040_0AF0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1125_1 ( .OUT(na1125_1), .IN1(1'b1), .IN2(~na377_1), .IN3(na375_1), .IN4(1'b1), .IN5(na161_1), .IN6(na1577_2), .IN7(na163_1),
                      .IN8(na162_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x25y94     80'h00_0018_00_0040_0AF0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1126_1 ( .OUT(na1126_1), .IN1(1'b1), .IN2(~na377_1), .IN3(~na375_1), .IN4(1'b1), .IN5(na165_2), .IN6(na143_1), .IN7(na145_1),
                      .IN8(na148_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x23y90     80'h00_0018_00_0040_0AF0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1127_1 ( .OUT(na1127_1), .IN1(1'b1), .IN2(~na377_1), .IN3(~na375_1), .IN4(1'b1), .IN5(na1576_2), .IN6(na150_1), .IN7(na146_2),
                      .IN8(na151_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x25y91     80'h00_0018_00_0040_0AF0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1128_1 ( .OUT(na1128_1), .IN1(1'b1), .IN2(~na377_1), .IN3(~na375_1), .IN4(1'b1), .IN5(na169_1), .IN6(na143_1), .IN7(na168_1),
                      .IN8(na148_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x23y89     80'h00_0018_00_0040_0AE0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1129_1 ( .OUT(na1129_1), .IN1(1'b1), .IN2(~na377_1), .IN3(~na375_1), .IN4(1'b1), .IN5(1'b0), .IN6(na144_2), .IN7(na147_2),
                      .IN8(na149_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x25y92     80'h00_0018_00_0040_0AF8_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1130_1 ( .OUT(na1130_1), .IN1(1'b1), .IN2(~na377_1), .IN3(~na375_1), .IN4(1'b1), .IN5(na172_1), .IN6(na1575_2), .IN7(na147_2),
                      .IN8(~na151_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x44y115     80'h00_0018_00_0040_0A70_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1131_1 ( .OUT(na1131_1), .IN1(1'b1), .IN2(~na184_1), .IN3(~na17_1), .IN4(1'b1), .IN5(na211_2), .IN6(na201_1), .IN7(na1598_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x34y118     80'h00_0018_00_0040_0AF4_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1132_1 ( .OUT(na1132_1), .IN1(1'b1), .IN2(~na184_1), .IN3(na17_1), .IN4(1'b1), .IN5(na202_2), .IN6(na181_1), .IN7(~na208_2),
                      .IN8(na193_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x44y117     80'h00_FE00_00_0040_0AF1_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1133_1 ( .OUT(na1133_1_i), .IN1(na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na19_1), .IN5(~na186_1), .IN6(na221_1), .IN7(na1131_1),
                      .IN8(na1132_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1133_2 ( .OUT(na1133_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1133_1_i) );
// C_MX4b////      x39y117     80'h00_0018_00_0040_0AF4_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1134_1 ( .OUT(na1134_1), .IN1(1'b1), .IN2(~na184_1), .IN3(~na17_1), .IN4(1'b1), .IN5(na1597_2), .IN6(na201_1), .IN7(~na216_1),
                      .IN8(na190_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x31y118     80'h00_0018_00_0040_0AF8_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1135_1 ( .OUT(na1135_1), .IN1(1'b1), .IN2(na184_1), .IN3(na17_1), .IN4(1'b1), .IN5(na202_2), .IN6(na181_1), .IN7(na1603_2),
                      .IN8(~na196_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x41y116     80'h00_FE00_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1136_1 ( .OUT(na1136_1_i), .IN1(na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(na19_1), .IN5(na1134_1), .IN6(na1135_1), .IN7(na191_1),
                      .IN8(na222_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1136_2 ( .OUT(na1136_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1136_1_i) );
// C_MX4b////      x36y117     80'h00_0018_00_0040_0A70_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1137_1 ( .OUT(na1137_1), .IN1(1'b1), .IN2(na184_1), .IN3(~na17_1), .IN4(1'b1), .IN5(na192_1), .IN6(na1586_2), .IN7(na1605_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x44y118     80'h00_FE00_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1138_1 ( .OUT(na1138_1_i), .IN1(na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na19_1), .IN5(na199_1), .IN6(na221_1), .IN7(na1137_1),
                      .IN8(na194_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1138_2 ( .OUT(na1138_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1138_1_i) );
// C_MX4b////      x35y117     80'h00_0018_00_0040_0AE2_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1139_1 ( .OUT(na1139_1), .IN1(1'b1), .IN2(~na184_1), .IN3(na17_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na200_1), .IN7(na176_2),
                      .IN8(na193_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x33y118     80'h00_0018_00_0040_0A74_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1140_1 ( .OUT(na1140_1), .IN1(1'b1), .IN2(~na184_1), .IN3(~na17_1), .IN4(1'b1), .IN5(na192_1), .IN6(na181_1), .IN7(~na1606_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x41y115     80'h00_FE00_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1141_1 ( .OUT(na1141_1_i), .IN1(na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(na19_1), .IN5(na1139_1), .IN6(na1140_1), .IN7(na223_2),
                      .IN8(na222_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1141_2 ( .OUT(na1141_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1141_1_i) );
// C_MX4b////      x35y115     80'h00_0018_00_0040_0AF8_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1142_1 ( .OUT(na1142_1), .IN1(1'b1), .IN2(~na184_1), .IN3(~na17_1), .IN4(1'b1), .IN5(na192_1), .IN6(na1600_2), .IN7(na1602_2),
                      .IN8(~na177_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x46y116     80'h00_FE00_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1143_1 ( .OUT(na1143_1_i), .IN1(~na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(na19_1), .IN5(na1142_1), .IN6(na204_1), .IN7(na209_2),
                      .IN8(na207_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1143_2 ( .OUT(na1143_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1143_1_i) );
// C_MX4b////      x29y113     80'h00_0018_00_0040_0AFE_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1144_1 ( .OUT(na1144_1), .IN1(1'b1), .IN2(~na184_1), .IN3(~na17_1), .IN4(1'b1), .IN5(na1589_2), .IN6(~na1601_2), .IN7(~na208_2),
                      .IN8(~na196_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x27y116     80'h00_0018_00_0040_0AFA_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1145_1 ( .OUT(na1145_1), .IN1(1'b1), .IN2(~na184_1), .IN3(~na17_1), .IN4(1'b1), .IN5(na192_1), .IN6(~na1601_2), .IN7(na1596_2),
                      .IN8(~na177_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x39y112     80'h00_FE00_00_0040_0AF8_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1146_1 ( .OUT(na1146_1_i), .IN1(na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(na19_1), .IN5(na1144_1), .IN6(na1145_1), .IN7(na223_2),
                      .IN8(~na210_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1146_2 ( .OUT(na1146_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1146_1_i) );
// C_MX4b/D///      x41y107     80'h00_FE00_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1147_1 ( .OUT(na1147_1_i), .IN1(na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na19_1), .IN5(na203_2), .IN6(na187_2), .IN7(na212_1),
                      .IN8(na213_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1147_2 ( .OUT(na1147_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1147_1_i) );
// C_MX4b////      x29y118     80'h00_0018_00_0040_0AF6_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1148_1 ( .OUT(na1148_1), .IN1(1'b1), .IN2(~na184_1), .IN3(na17_1), .IN4(1'b1), .IN5(na192_1), .IN6(~na1587_2), .IN7(~na198_1),
                      .IN8(na215_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x31y115     80'h00_0018_00_0040_0AF9_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1149_1 ( .OUT(na1149_1), .IN1(1'b1), .IN2(na184_1), .IN3(na17_1), .IN4(1'b1), .IN5(~na217_2), .IN6(na181_1), .IN7(na1590_2),
                      .IN8(~na177_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x39y109     80'h00_FE00_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1150_1 ( .OUT(na1150_1_i), .IN1(~na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(na19_1), .IN5(na1149_1), .IN6(na1148_1), .IN7(na188_2),
                      .IN8(na214_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1150_2 ( .OUT(na1150_1), .CLK(na1197_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1150_1_i) );
// C_MX4b////      x35y110     80'h00_0018_00_0040_0A50_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1151_1 ( .OUT(na1151_1), .IN1(~na8_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1_2), .IN5(na774_1), .IN6(1'b0), .IN7(na1675_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x35y108     80'h00_0018_00_0040_0A55_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1152_1 ( .OUT(na1152_1), .IN1(~na8_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1_2), .IN5(~na1612_2), .IN6(1'b0), .IN7(~na241_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x31y105     80'h00_0018_00_0040_0A90_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1153_1 ( .OUT(na1153_1), .IN1(~na1614_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1640_2), .IN5(na297_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(na1609_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x27y104     80'h00_0018_00_0040_0AB0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1154_1 ( .OUT(na1154_1), .IN1(~na22_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na292_1), .IN5(na556_2), .IN6(na253_1), .IN7(1'b0),
                      .IN8(na252_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x31y112     80'h00_0018_00_0040_0AA0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1155_1 ( .OUT(na1155_1), .IN1(na8_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1_2), .IN5(1'b0), .IN6(na776_2), .IN7(1'b0), .IN8(na1680_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x31y114     80'h00_0018_00_0040_0AA0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1156_1 ( .OUT(na1156_1), .IN1(na8_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1_2), .IN5(1'b0), .IN6(na776_1), .IN7(1'b0), .IN8(na1678_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x33y114     80'h00_0018_00_0040_0A50_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1157_1 ( .OUT(na1157_1), .IN1(~na8_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1_2), .IN5(na774_2), .IN6(1'b0), .IN7(na1676_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x25y104     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1158_1 ( .OUT(na1158_1), .IN1(na22_1), .IN2(1'b1), .IN3(1'b1), .IN4(na292_1), .IN5(na332_2), .IN6(na333_2), .IN7(na334_1),
                      .IN8(na560_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x25y102     80'h00_0018_00_0040_0AE0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1159_1 ( .OUT(na1159_1), .IN1(~na22_1), .IN2(1'b1), .IN3(1'b1), .IN4(na292_1), .IN5(1'b0), .IN6(na339_1), .IN7(na559_1),
                      .IN8(na340_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x27y102     80'h00_0018_00_0040_0AD0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1160_1 ( .OUT(na1160_1), .IN1(na22_1), .IN2(1'b1), .IN3(1'b1), .IN4(na292_1), .IN5(na345_1), .IN6(1'b0), .IN7(na346_2), .IN8(na558_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x25y100     80'h00_0018_00_0040_0AB0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1161_1 ( .OUT(na1161_1), .IN1(~na22_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na292_1), .IN5(na557_1), .IN6(na350_2), .IN7(1'b0),
                      .IN8(na349_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x32y103     80'h00_0018_00_0040_0AE0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1162_1 ( .OUT(na1162_1), .IN1(~na22_1), .IN2(1'b1), .IN3(1'b1), .IN4(na292_1), .IN5(1'b0), .IN6(na357_1), .IN7(na555_2),
                      .IN8(na358_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x28y102     80'h00_0018_00_0040_0AD0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1163_1 ( .OUT(na1163_1), .IN1(na22_1), .IN2(1'b1), .IN3(1'b1), .IN4(na292_1), .IN5(na363_2), .IN6(1'b0), .IN7(na364_1), .IN8(na554_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y91     80'h00_0018_00_0040_0A60_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1164_1 ( .OUT(na1164_1), .IN1(1'b1), .IN2(na448_2), .IN3(1'b1), .IN4(~na1649_2), .IN5(1'b0), .IN6(na337_2), .IN7(na324_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x43y105     80'h00_0018_00_0040_0A50_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1165_1 ( .OUT(na1165_1), .IN1(1'b1), .IN2(na29_1), .IN3(na25_1), .IN4(1'b1), .IN5(na689_1), .IN6(1'b0), .IN7(na1665_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x39y97     80'h00_0018_00_0040_0A50_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1166_1 ( .OUT(na1166_1), .IN1(1'b1), .IN2(na29_1), .IN3(na25_1), .IN4(1'b1), .IN5(na685_2), .IN6(1'b0), .IN7(na1661_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x33y103     80'h00_0018_00_0040_0AA0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1167_1 ( .OUT(na1167_1), .IN1(1'b1), .IN2(~na29_1), .IN3(na25_1), .IN4(1'b1), .IN5(1'b0), .IN6(na687_2), .IN7(1'b0), .IN8(na1664_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x35y105     80'h00_0018_00_0040_0AA0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1168_1 ( .OUT(na1168_1), .IN1(1'b1), .IN2(~na29_1), .IN3(na25_1), .IN4(1'b1), .IN5(1'b0), .IN6(na687_1), .IN7(1'b0), .IN8(na1663_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x37y95     80'h00_0018_00_0040_0A50_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1169_1 ( .OUT(na1169_1), .IN1(1'b1), .IN2(na29_1), .IN3(na25_1), .IN4(1'b1), .IN5(na685_1), .IN6(1'b0), .IN7(na1659_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x41y95     80'h00_0018_00_0040_0AAA_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1170_1 ( .OUT(na1170_1), .IN1(1'b1), .IN2(~na29_1), .IN3(na25_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1645_2), .IN7(1'b0), .IN8(~na416_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x41y90     80'h00_0018_00_0040_0AD0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1171_1 ( .OUT(na1171_1), .IN1(na31_1), .IN2(1'b1), .IN3(1'b1), .IN4(na420_2), .IN5(na449_1), .IN6(1'b0), .IN7(na450_2), .IN8(na552_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x44y92     80'h00_0018_00_0040_0AE0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1172_1 ( .OUT(na1172_1), .IN1(~na31_1), .IN2(1'b1), .IN3(1'b1), .IN4(na420_2), .IN5(1'b0), .IN6(na471_1), .IN7(na547_2),
                      .IN8(na472_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x44y91     80'h00_0018_00_0040_0AD0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1173_1 ( .OUT(na1173_1), .IN1(na31_1), .IN2(1'b1), .IN3(1'b1), .IN4(na420_2), .IN5(na475_2), .IN6(1'b0), .IN7(na476_1), .IN8(na548_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y89     80'h00_0018_00_0040_0AD0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1174_1 ( .OUT(na1174_1), .IN1(na31_1), .IN2(1'b1), .IN3(1'b1), .IN4(na420_2), .IN5(na479_1), .IN6(1'b0), .IN7(na480_1), .IN8(na549_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x41y91     80'h00_0018_00_0040_0A70_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1175_1 ( .OUT(na1175_1), .IN1(na31_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na420_2), .IN5(na484_1), .IN6(na550_1), .IN7(na483_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y95     80'h00_0018_00_0040_0A70_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1176_1 ( .OUT(na1176_1), .IN1(na31_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na420_2), .IN5(na488_1), .IN6(na551_1), .IN7(na487_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y92     80'h00_0018_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1177_1 ( .OUT(na1177_1), .IN1(na31_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na420_2), .IN5(na493_2), .IN6(na553_2), .IN7(na491_1),
                      .IN8(na492_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000050)) 
           _a1178 ( .Y(na1178_1), .I(btn) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a1179 ( .Y(na1179_1), .I(clk) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1180 ( .O(led), .A(na1539_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1181 ( .O(oled_clk), .A(na1540_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1182 ( .O(oled_clk_1), .A(na1541_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1183 ( .O(oled_csn), .A(na1542_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1184 ( .O(oled_dc), .A(na1543_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1185 ( .O(oled_dc_1), .A(na1544_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1186 ( .O(oled_mosi), .A(na1545_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1187 ( .O(oled_mosi_1), .A(na1546_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1188 ( .O(oled_resn), .A(na1547_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1189 ( .O(oled_resn_1), .A(na1548_10) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_07_08_0A_1C_82)) 
           _a1192 ( .USR_PLL_LOCKED_STDY(_d0), .USR_PLL_LOCKED(_d1), .CLK270(na1192_3), .CLK180(na1192_4), .CLK90(na1192_5), .CLK0(na1192_6),
                    .CLK_REF_OUT(_d2), .CLK_REF(na1201_1), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
// C_AND////      x37y106     80'h00_0018_00_0000_0888_8844
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1193_1 ( .OUT(na1193_1), .IN1(~na1199_1), .IN2(na1194_1), .IN3(~na1196_1), .IN4(na7_1), .IN5(na1195_2), .IN6(na1194_2), .IN7(na1200_1),
                      .IN8(na1198_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x33y102     80'h00_0078_00_0000_0C66_3C5C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1194_1 ( .OUT(na1194_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na782_2), .IN7(1'b0), .IN8(~na270_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1194_4 ( .OUT(na1194_2), .IN1(1'b0), .IN2(na782_1), .IN3(~na272_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x39y99     80'h00_0060_00_0000_0C0E_FF0D
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1195_4 ( .OUT(na1195_2), .IN1(~na780_1), .IN2(na219_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x38y103     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1196_1 ( .OUT(na1196_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na780_2), .IN6(1'b1), .IN7(1'b1), .IN8(na270_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0011_0014)) 
           _a1197 ( .GLB0(na1197_1), .GLB1(na1197_2), .GLB2(_d3), .GLB3(_d4), .CLK_FB0(_d5), .CLK_FB1(_d6), .CLK_FB2(_d7), .CLK_FB3(_d8),
                    .CLK0_0(na1192_6), .CLK0_90(na1192_5), .CLK0_180(na1192_4), .CLK0_270(na1192_3), .CLK0_BYP(1'b0), .CLK1_0(1'b0),
                    .CLK1_90(1'b0), .CLK1_180(1'b0), .CLK1_270(1'b0), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0),
                    .CLK2_270(1'b0), .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0),
                    .USR_GLB0(1'b0), .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0),
                    .USR_FB3(1'b0) );
// C_///OR/      x40y102     80'h00_0060_00_0000_0C0E_FF0B
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1198_4 ( .OUT(na1198_2), .IN1(na785_1), .IN2(~na219_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y103     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1199_1 ( .OUT(na1199_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na780_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na270_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x36y103     80'h00_0018_00_0000_0C66_5300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1200_1 ( .OUT(na1200_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1116_2), .IN7(~na241_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a1201 ( .PCLK0(na1201_1), .PCLK1(_d9), .PCLK2(_d10), .PCLK3(_d11), .CLK0(na1179_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0),
                    .SER_CLK(1'b0), .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_OR////      x44y107     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1203_1 ( .OUT(na1203_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na681_2), .IN7(1'b0), .IN8(~na13_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x40y112     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1204_4 ( .OUT(na1204_2), .IN1(~na265_1), .IN2(1'b1), .IN3(na17_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x44y111     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1205_4 ( .OUT(na1205_2), .IN1(~na683_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na13_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x44y112     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1206_1 ( .OUT(na1206_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na265_1), .IN6(1'b1), .IN7(1'b1), .IN8(na19_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x34y103     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1207_2 ( .OUT(na1207_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1207_6 ( .COUTY1(na1207_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1207_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x40y107     80'h00_0078_00_0000_0C66_A55A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1208_1 ( .OUT(na1208_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na402_1), .IN6(1'b0), .IN7(na696_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1208_4 ( .OUT(na1208_2), .IN1(na402_2), .IN2(1'b0), .IN3(~na691_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x39y99     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1209_1 ( .OUT(na1209_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na994_2), .IN6(1'b0), .IN7(1'b0), .IN8(na416_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x41y108     80'h00_0078_00_0000_0C66_C3C5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1210_1 ( .OUT(na1210_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na410_1), .IN7(1'b0), .IN8(na693_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1210_4 ( .OUT(na1210_2), .IN1(~na412_1), .IN2(1'b0), .IN3(1'b0), .IN4(na693_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x39y107     80'h00_0018_00_0000_0C66_A500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1212_1 ( .OUT(na1212_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na412_2), .IN6(1'b0), .IN7(na691_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y108     80'h00_0018_00_0040_0A31_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1214_1 ( .OUT(na1214_1), .IN1(~na39_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na35_1), .IN6(na219_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x31y101     80'h00_0018_00_0000_0EEE_EEBE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1217_1 ( .OUT(na1217_1), .IN1(na170_1), .IN2(na171_1), .IN3(na167_1), .IN4(~na1218_2), .IN5(na166_1), .IN6(na160_1), .IN7(na167_2),
                      .IN8(na164_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x32y108     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1218_4 ( .OUT(na1218_2), .IN1(1'b1), .IN2(~na173_2), .IN3(na241_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x26y93     80'h00_0018_00_0000_0888_4245
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1219_1 ( .OUT(na1219_1), .IN1(~na258_1), .IN2(1'b1), .IN3(~na375_2), .IN4(na139_2), .IN5(na137_2), .IN6(~na377_2), .IN7(~na141_2),
                      .IN8(na155_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x43y87     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1220_1 ( .OUT(na1220_1), .IN1(1'b1), .IN2(na48_2), .IN3(1'b0), .IN4(1'b0), .IN5(na135_2), .IN6(na48_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x33y92     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1221_1 ( .OUT(na1221_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na58_1), .IN6(na51_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x32y91     80'h00_0018_00_0000_0C88_21FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1224_1 ( .OUT(na1224_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na166_1), .IN6(~na1225_2), .IN7(na167_1),
                      .IN8(~na1581_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y90     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1225_4 ( .OUT(na1225_2), .IN1(1'b1), .IN2(1'b1), .IN3(na167_2), .IN4(na164_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y95     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1226_1 ( .OUT(na1226_1), .IN1(1'b1), .IN2(na1563_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na63_2), .IN8(~na61_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x38y98     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1227_4 ( .OUT(na1227_2), .IN1(1'b1), .IN2(1'b1), .IN3(na167_1), .IN4(na62_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y89     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1228_4 ( .OUT(na1228_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na167_2), .IN4(~na164_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x41y93     80'h00_0018_00_0040_0A51_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1229_1 ( .OUT(na1229_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na96_2), .IN5(~na64_1), .IN6(1'b0), .IN7(na63_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x32y98     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1230_4 ( .OUT(na1230_2), .IN1(~na166_1), .IN2(~na1225_2), .IN3(na167_1), .IN4(na1581_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y102     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1232_1 ( .OUT(na1232_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na72_1), .IN8(na66_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x43y100     80'h00_0018_00_0000_0C88_54FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1234_1 ( .OUT(na1234_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na69_2), .IN6(na1441_2), .IN7(~na14_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x52y113     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1236_1 ( .OUT(na1236_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na73_1), .IN7(1'b1), .IN8(~na1143_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x49y113     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1237_4 ( .OUT(na1237_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1133_1), .IN4(na1138_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y88     80'h00_0018_00_0040_0A51_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1238_1 ( .OUT(na1238_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na96_2), .IN5(~na75_1), .IN6(1'b0), .IN7(na74_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x34y89     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1239_1 ( .OUT(na1239_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na166_1), .IN6(~na1225_2), .IN7(~na167_1),
                      .IN8(~na1581_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y87     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1240_1 ( .OUT(na1240_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na77_1), .IN6(na78_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x34y92     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1241_1 ( .OUT(na1241_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na167_1), .IN8(na62_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y88     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1242_1 ( .OUT(na1242_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na79_1), .IN6(na78_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x32y90     80'h00_0060_00_0000_0C08_FF41
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1243_4 ( .OUT(na1243_2), .IN1(~na166_1), .IN2(~na1225_2), .IN3(~na167_1), .IN4(na1581_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y99     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1244_1 ( .OUT(na1244_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na80_1), .IN8(~na81_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y114     80'h00_0018_00_0000_0C88_14FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1245_1 ( .OUT(na1245_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1141_1), .IN6(na1136_1), .IN7(~na1246_1),
                      .IN8(~na1143_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y115     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1246_1 ( .OUT(na1246_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1133_1), .IN8(na1138_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y89     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1247_1 ( .OUT(na1247_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na84_1), .IN8(na83_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x32y89     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1248_4 ( .OUT(na1248_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na167_1), .IN4(~na85_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x39y90     80'h00_0018_00_0040_0AA2_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1250_1 ( .OUT(na1250_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na96_2), .IN5(1'b0), .IN6(~na87_1), .IN7(1'b0), .IN8(na89_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x34y92     80'h00_0060_00_0000_0C08_FF53
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1251_4 ( .OUT(na1251_2), .IN1(1'b1), .IN2(~na88_1), .IN3(~na167_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x30y93     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1252_4 ( .OUT(na1252_2), .IN1(1'b1), .IN2(~na160_1), .IN3(na167_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x27y90     80'h00_0060_00_0000_0C06_FFA3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1253_4 ( .OUT(na1253_2), .IN1(1'b0), .IN2(~na160_1), .IN3(na167_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x39y91     80'h00_0018_00_0040_0AA2_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1254_1 ( .OUT(na1254_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na96_2), .IN5(1'b0), .IN6(~na90_1), .IN7(1'b0), .IN8(na89_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x31y91     80'h00_0060_00_0000_0C08_FF4C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1255_4 ( .OUT(na1255_2), .IN1(1'b1), .IN2(na160_1), .IN3(~na167_1), .IN4(na1256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x30y96     80'h00_0018_00_0040_0C64_3500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1256_1 ( .OUT(na1256_1), .IN1(1'b0), .IN2(1'b1), .IN3(~na167_2), .IN4(1'b0), .IN5(~na166_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na164_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y93     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1257_1 ( .OUT(na1257_1), .IN1(1'b1), .IN2(na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(na92_2), .IN6(~na93_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x35y96     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1258_4 ( .OUT(na1258_2), .IN1(1'b1), .IN2(na94_1), .IN3(~na167_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x30y95     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1260_4 ( .OUT(na1260_2), .IN1(1'b1), .IN2(na160_1), .IN3(na167_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x43y96     80'h00_0018_00_0040_0AA8_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1261_1 ( .OUT(na1261_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na96_2), .IN5(1'b0), .IN6(na95_1), .IN7(1'b0), .IN8(~na96_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y94     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1264_1 ( .OUT(na1264_1), .IN1(1'b1), .IN2(na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(na99_2), .IN6(~na100_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x32y92     80'h00_0018_00_0040_0C98_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1266_1 ( .OUT(na1266_1), .IN1(1'b1), .IN2(1'b0), .IN3(1'b0), .IN4(~na164_1), .IN5(1'b1), .IN6(na160_1), .IN7(~na167_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y91     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1267_1 ( .OUT(na1267_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na103_1), .IN8(na102_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x39y87     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1270_1 ( .OUT(na1270_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na106_1), .IN8(na131_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y94     80'h00_0018_00_0000_0888_A513
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1271_1 ( .OUT(na1271_1), .IN1(1'b1), .IN2(~na160_1), .IN3(~na167_1), .IN4(~na164_1), .IN5(~na166_1), .IN6(1'b1), .IN7(na167_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y100     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1272_1 ( .OUT(na1272_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na80_2), .IN8(~na109_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x50y114     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1273_4 ( .OUT(na1273_2), .IN1(1'b1), .IN2(na110_1), .IN3(1'b1), .IN4(~na1143_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x48y115     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1274_4 ( .OUT(na1274_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1133_1), .IN4(~na1138_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y100     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1275_1 ( .OUT(na1275_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na112_1), .IN8(na111_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x48y113     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1276_4 ( .OUT(na1276_2), .IN1(~na1141_1), .IN2(~na1136_1), .IN3(~na1246_1), .IN4(~na1143_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y97     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1278_1 ( .OUT(na1278_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na115_1), .IN6(na578_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x32y94     80'h00_0018_00_0040_0A81_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1280_1 ( .OUT(na1280_1), .IN1(1'b1), .IN2(~na160_1), .IN3(~na167_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b0), .IN7(1'b0), .IN8(na164_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x34y96     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1281_1 ( .OUT(na1281_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na118_1), .IN6(na117_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x27y97     80'h00_0018_00_0000_0C88_C2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1282_1 ( .OUT(na1282_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na166_1), .IN6(~na1253_2), .IN7(1'b1), .IN8(na164_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x38y96     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1284_1 ( .OUT(na1284_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na122_1), .IN8(na121_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y94     80'h00_0018_00_0000_0C88_C8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1285_1 ( .OUT(na1285_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na166_1), .IN6(na160_1), .IN7(1'b1), .IN8(na164_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y93     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1286_1 ( .OUT(na1286_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na127_1), .IN6(na51_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y87     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1289_1 ( .OUT(na1289_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na132_1), .IN8(na131_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x30y94     80'h00_0018_00_0000_0888_541F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1290_1 ( .OUT(na1290_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na167_2), .IN4(~na164_1), .IN5(~na166_1), .IN6(na160_1), .IN7(~na167_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x38y88     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1291_1 ( .OUT(na1291_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na134_1), .IN6(na133_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x30y89     80'h00_0018_00_0000_0C88_14FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1292_1 ( .OUT(na1292_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na166_1), .IN6(na1253_2), .IN7(~na167_1),
                      .IN8(~na164_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x44y88     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1293_1 ( .OUT(na1293_1), .IN1(1'b1), .IN2(na48_2), .IN3(1'b0), .IN4(1'b0), .IN5(na135_1), .IN6(na136_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x30y85     80'h00_0018_00_0040_0A71_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1298_1 ( .OUT(na1298_1), .IN1(1'b1), .IN2(na1565_2), .IN3(1'b1), .IN4(na138_2), .IN5(~na1571_2), .IN6(na1572_2), .IN7(na142_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x30y86     80'h00_0018_00_0040_0ADB_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1299_1 ( .OUT(na1299_1), .IN1(1'b1), .IN2(na1565_2), .IN3(1'b1), .IN4(na138_2), .IN5(~na1571_2), .IN6(1'b1), .IN7(na142_1),
                      .IN8(~na1573_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x29y85     80'h00_0018_00_0040_0ADB_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1300_1 ( .OUT(na1300_1), .IN1(1'b1), .IN2(na1566_2), .IN3(1'b1), .IN4(na138_1), .IN5(~na1571_2), .IN6(1'b1), .IN7(na142_1),
                      .IN8(~na1573_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x27y87     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1301_4 ( .OUT(na1301_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na142_1), .IN4(na138_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x21y94     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1302_1 ( .OUT(na1302_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na57_2), .IN7(~na772_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x27y97     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1303_4 ( .OUT(na1303_2), .IN1(1'b1), .IN2(~na256_1), .IN3(1'b1), .IN4(na155_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x27y86     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1304_1 ( .OUT(na1304_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1565_2), .IN7(1'b1), .IN8(na138_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x32y88     80'h00_0018_00_0040_0C64_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1308_1 ( .OUT(na1308_1), .IN1(1'b0), .IN2(1'b1), .IN3(~na142_1), .IN4(1'b0), .IN5(1'b1), .IN6(na1566_2), .IN7(1'b1), .IN8(na138_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x27y88     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1311_4 ( .OUT(na1311_2), .IN1(1'b1), .IN2(na1565_2), .IN3(1'b1), .IN4(~na138_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x29y86     80'h00_0018_00_0040_0AB2_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1312_1 ( .OUT(na1312_1), .IN1(1'b1), .IN2(~na1566_2), .IN3(na142_1), .IN4(1'b1), .IN5(na1564_2), .IN6(~na1565_2), .IN7(1'b0),
                      .IN8(na138_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x32y97     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1313_1 ( .OUT(na1313_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na175_1), .IN6(na227_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x34y98     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1314_4 ( .OUT(na1314_2), .IN1(1'b1), .IN2(~na88_1), .IN3(na167_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y111     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1321_1 ( .OUT(na1321_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na180_1), .IN8(na178_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x39y114     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1325_1 ( .OUT(na1325_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na187_2), .IN7(1'b1), .IN8(~na195_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x36y113     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1327_4 ( .OUT(na1327_2), .IN1(~na189_2), .IN2(1'b1), .IN3(~na180_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x40y113     80'h00_0018_00_0000_0888_CFA6
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1329_1 ( .OUT(na1329_1), .IN1(~na189_2), .IN2(na206_1), .IN3(~na179_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(~na178_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x38y113     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1333_1 ( .OUT(na1333_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na189_2), .IN6(1'b1), .IN7(~na180_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y116     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1334_1 ( .OUT(na1334_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na189_2), .IN6(1'b1), .IN7(na180_1), .IN8(na178_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x39y113     80'h00_0018_00_0000_0CEE_A700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1335_1 ( .OUT(na1335_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1552_2), .IN6(~na206_1), .IN7(na180_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y107     80'h00_0018_00_0040_0A31_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1340_1 ( .OUT(na1340_1), .IN1(~na39_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na220_2), .IN6(na219_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y90     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1345_1 ( .OUT(na1345_1), .IN1(1'b1), .IN2(na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(na224_1), .IN6(~na225_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x34y89     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1346_4 ( .OUT(na1346_2), .IN1(1'b1), .IN2(na226_1), .IN3(~na167_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x30y90     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1347_4 ( .OUT(na1347_2), .IN1(1'b1), .IN2(~na160_1), .IN3(1'b1), .IN4(na164_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x31y98     80'h00_0018_00_0040_0AA8_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1348_1 ( .OUT(na1348_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na96_2), .IN5(1'b0), .IN6(na227_1), .IN7(1'b0), .IN8(~na228_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x31y99     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1349_4 ( .OUT(na1349_2), .IN1(1'b1), .IN2(na160_1), .IN3(na167_1), .IN4(na1256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x33y89     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1350_1 ( .OUT(na1350_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na230_1), .IN6(na229_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y91     80'h00_0018_00_0000_0888_5513
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1351_1 ( .OUT(na1351_1), .IN1(1'b1), .IN2(~na160_1), .IN3(~na167_1), .IN4(~na164_1), .IN5(~na166_1), .IN6(1'b1), .IN7(~na167_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x24y111     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1352_4 ( .OUT(na1352_2), .IN1(~na238_1), .IN2(1'b1), .IN3(1'b1), .IN4(na786_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x28y104     80'h00_0018_00_0040_0AC8_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1353_1 ( .OUT(na1353_1), .IN1(na39_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na241_1), .IN8(~na242_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x21y91     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1356_1 ( .OUT(na1356_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na764_1), .IN8(na323_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x21y95     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1357_1 ( .OUT(na1357_1), .IN1(1'b1), .IN2(na366_2), .IN3(1'b0), .IN4(1'b0), .IN5(na244_2), .IN6(~na247_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x30y97     80'h00_0018_00_0000_0888_4F34
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1358_1 ( .OUT(na1358_1), .IN1(~na23_1), .IN2(na1359_2), .IN3(1'b1), .IN4(~na1_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na276_1),
                      .IN8(na292_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x25y98     80'h00_0078_00_0000_0C88_F211
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1359_1 ( .OUT(na1359_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na249_1), .IN6(~na248_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1359_4 ( .OUT(na1359_2), .IN1(~na328_2), .IN2(~na1631_2), .IN3(~na322_1), .IN4(~na323_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x27y100     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1360_1 ( .OUT(na1360_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na250_2), .IN8(na929_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x25y101     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1361_1 ( .OUT(na1361_1), .IN1(1'b1), .IN2(na366_2), .IN3(1'b0), .IN4(1'b0), .IN5(na254_2), .IN6(~na255_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x29y97     80'h00_0078_00_0000_0C88_AC4C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1363_1 ( .OUT(na1363_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na94_1), .IN7(na167_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1363_4 ( .OUT(na1363_2), .IN1(1'b1), .IN2(na1359_2), .IN3(~na1219_1), .IN4(na1615_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x27y95     80'h00_0018_00_0040_0A31_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1364_1 ( .OUT(na1364_1), .IN1(~na262_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na262_1), .IN6(na260_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x36y110     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1365_1 ( .OUT(na1365_1), .IN1(~na23_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na241_1), .IN8(~na1_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x39y96     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1366_1 ( .OUT(na1366_1), .IN1(1'b1), .IN2(na1563_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na263_1), .IN8(~na264_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x31y96     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1367_1 ( .OUT(na1367_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na167_1), .IN8(~na85_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x42y116     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1370_1 ( .OUT(na1370_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1136_1), .IN7(na1133_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x45y115     80'h00_0018_00_0000_0C66_AC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1371_1 ( .OUT(na1371_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1136_1), .IN7(na1133_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y107     80'h00_0018_00_0040_0AC4_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1372_1 ( .OUT(na1372_1), .IN1(~na39_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na271_1), .IN8(na270_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x31y109     80'h00_0018_00_0040_0AC8_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1375_1 ( .OUT(na1375_1), .IN1(na39_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na272_2), .IN8(~na273_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y96     80'h00_0018_00_0040_0A51_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1378_1 ( .OUT(na1378_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na96_2), .IN5(~na275_1), .IN6(1'b0), .IN7(na263_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x32y95     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1379_1 ( .OUT(na1379_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na226_1), .IN7(na167_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x35y103     80'h00_0060_00_0000_0C0E_FF57
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1380_4 ( .OUT(na1380_2), .IN1(~na39_2), .IN2(~na173_2), .IN3(~na250_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x33y106     80'h00_0060_00_0000_0C08_FFA7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1381_4 ( .OUT(na1381_2), .IN1(~na39_2), .IN2(~na1382_1), .IN3(na276_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x33y110     80'h00_0018_00_0040_0AC8_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1382_1 ( .OUT(na1382_1), .IN1(~na23_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na241_1), .IN8(~na1_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y104     80'h00_0018_00_0040_0AC4_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1383_1 ( .OUT(na1383_1), .IN1(~na39_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na281_1), .IN8(na270_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y105     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1386_1 ( .OUT(na1386_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na282_2), .IN8(~na283_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y117     80'h00_0018_00_0000_0888_344F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1387_1 ( .OUT(na1387_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1133_1), .IN4(na1143_1), .IN5(~na1141_1), .IN6(na1136_1), .IN7(1'b1),
                      .IN8(~na1138_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y101     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1388_1 ( .OUT(na1388_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1619_2), .IN6(na287_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x25y112     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1408_1 ( .OUT(na1408_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na238_1), .IN6(1'b1), .IN7(na792_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x27y111     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1409_4 ( .OUT(na1409_2), .IN1(~na238_1), .IN2(1'b1), .IN3(1'b1), .IN4(na790_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x20y109     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1410_1 ( .OUT(na1410_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na238_1), .IN6(1'b1), .IN7(1'b1), .IN8(na790_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y88     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1411_1 ( .OUT(na1411_1), .IN1(~na311_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1630_2), .IN8(na309_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x32y116     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1412_4 ( .OUT(na1412_2), .IN1(~na238_1), .IN2(1'b1), .IN3(na788_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x23y109     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1413_4 ( .OUT(na1413_2), .IN1(~na238_1), .IN2(1'b1), .IN3(na788_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x24y111     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1414_1 ( .OUT(na1414_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na238_1), .IN6(1'b1), .IN7(1'b1), .IN8(na786_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x30y106     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1415_4 ( .OUT(na1415_2), .IN1(~na238_1), .IN2(1'b1), .IN3(~na314_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x20y96     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1416_1 ( .OUT(na1416_1), .IN1(1'b1), .IN2(na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na322_1), .IN8(na766_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x21y93     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1417_1 ( .OUT(na1417_1), .IN1(1'b1), .IN2(~na57_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na764_2), .IN8(na323_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x48y87     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1418_1 ( .OUT(na1418_1), .IN1(na311_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na324_2), .IN8(na325_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x48y85     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1419_1 ( .OUT(na1419_1), .IN1(1'b1), .IN2(~na48_2), .IN3(1'b0), .IN4(1'b0), .IN5(na703_2), .IN6(na337_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x42y86     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1422_1 ( .OUT(na1422_1), .IN1(1'b1), .IN2(~na48_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na330_2), .IN8(na343_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x21y99     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1424_1 ( .OUT(na1424_1), .IN1(1'b1), .IN2(~na366_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na336_1), .IN8(na335_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y87     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1425_1 ( .OUT(na1425_1), .IN1(1'b1), .IN2(~na48_2), .IN3(1'b0), .IN4(1'b0), .IN5(na338_2), .IN6(na337_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x24y100     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1426_1 ( .OUT(na1426_1), .IN1(1'b1), .IN2(na366_2), .IN3(1'b0), .IN4(1'b0), .IN5(na341_1), .IN6(~na342_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x42y87     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1427_1 ( .OUT(na1427_1), .IN1(1'b1), .IN2(~na48_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na344_2), .IN8(na343_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x21y96     80'h00_0018_00_0040_0A54_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1428_1 ( .OUT(na1428_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1637_2), .IN5(na347_1), .IN6(1'b0), .IN7(~na348_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x23y100     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1429_1 ( .OUT(na1429_1), .IN1(1'b1), .IN2(na366_2), .IN3(1'b0), .IN4(1'b0), .IN5(na351_1), .IN6(~na352_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y87     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1430_1 ( .OUT(na1430_1), .IN1(na311_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na353_1), .IN6(na354_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y87     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1431_1 ( .OUT(na1431_1), .IN1(~na311_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na356_2), .IN6(na355_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x26y98     80'h00_0018_00_0040_0A54_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1432_1 ( .OUT(na1432_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1637_2), .IN5(na359_2), .IN6(1'b0), .IN7(~na360_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x51y86     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1433_1 ( .OUT(na1433_1), .IN1(na311_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na353_2), .IN6(na362_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x24y99     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1434_1 ( .OUT(na1434_1), .IN1(1'b1), .IN2(~na366_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1636_2), .IN8(na365_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x42y98     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1435_1 ( .OUT(na1435_1), .IN1(1'b1), .IN2(~na1550_2), .IN3(1'b0), .IN4(1'b0), .IN5(na675_2), .IN6(na1638_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x23y98     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1436_1 ( .OUT(na1436_1), .IN1(1'b1), .IN2(na369_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na368_1), .IN8(~na370_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x29y101     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1437_1 ( .OUT(na1437_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1363_2), .IN6(na371_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x44y97     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1438_1 ( .OUT(na1438_1), .IN1(1'b1), .IN2(na1550_2), .IN3(1'b0), .IN4(1'b0), .IN5(na372_1), .IN6(na677_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y88     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1439_1 ( .OUT(na1439_1), .IN1(~na311_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na374_2), .IN8(na309_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y93     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1440_1 ( .OUT(na1440_1), .IN1(1'b1), .IN2(na384_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na379_2), .IN8(~na380_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x47y96     80'h00_0078_00_0000_0C88_C511
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1441_1 ( .OUT(na1441_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na381_1), .IN6(1'b1), .IN7(1'b1), .IN8(na382_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1441_4 ( .OUT(na1441_2), .IN1(~na372_1), .IN2(~na1639_2), .IN3(~na331_1), .IN4(~na367_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x42y90     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1442_1 ( .OUT(na1442_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na383_1), .IN6(na1038_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y99     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1444_1 ( .OUT(na1444_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na385_2), .IN6(~na386_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x50y115     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1445_4 ( .OUT(na1445_2), .IN1(~na1371_1), .IN2(~na1700_2), .IN3(~na1698_2), .IN4(~na1138_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y109     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1447_1 ( .OUT(na1447_1), .IN1(1'b1), .IN2(~na389_2), .IN3(1'b0), .IN4(1'b0), .IN5(na390_1), .IN6(na388_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x43y95     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1448_1 ( .OUT(na1448_1), .IN1(1'b1), .IN2(na32_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na25_1), .IN8(na416_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x46y97     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1449_1 ( .OUT(na1449_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na391_1), .IN6(~na392_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x44y114     80'h00_0018_00_0000_0888_341F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1450_1 ( .OUT(na1450_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1133_1), .IN4(~na1143_1), .IN5(~na1141_1), .IN6(na1136_1), .IN7(1'b1),
                      .IN8(~na1138_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y99     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1451_1 ( .OUT(na1451_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na391_2), .IN6(~na394_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x42y114     80'h00_0018_00_0000_0888_2533
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1452_1 ( .OUT(na1452_1), .IN1(1'b1), .IN2(~na1136_1), .IN3(1'b1), .IN4(~na1143_1), .IN5(~na1141_1), .IN6(1'b1), .IN7(na1133_1),
                      .IN8(~na1138_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x44y98     80'h00_0018_00_0000_0888_FA7C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1455_1 ( .OUT(na1455_1), .IN1(1'b0), .IN2(na470_2), .IN3(~na1456_1), .IN4(~na1642_2), .IN5(na397_2), .IN6(1'b0), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x46y95     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1456_1 ( .OUT(na1456_1), .IN1(1'b1), .IN2(na32_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na25_1), .IN8(na416_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x43y93     80'h00_0018_00_0040_0A54_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1457_1 ( .OUT(na1457_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1642_2), .IN5(na402_1), .IN6(1'b0), .IN7(~na403_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x43y92     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1460_1 ( .OUT(na1460_1), .IN1(1'b1), .IN2(na399_2), .IN3(1'b0), .IN4(1'b0), .IN5(na412_2), .IN6(~na409_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x42y94     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1463_1 ( .OUT(na1463_1), .IN1(1'b1), .IN2(~na399_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na411_1), .IN6(na410_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x43y91     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1466_1 ( .OUT(na1466_1), .IN1(1'b1), .IN2(na399_2), .IN3(1'b0), .IN4(1'b0), .IN5(na412_1), .IN6(~na413_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x42y93     80'h00_0018_00_0040_0A54_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1469_1 ( .OUT(na1469_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1642_2), .IN5(na402_2), .IN6(1'b0), .IN7(~na415_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x44y94     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1472_1 ( .OUT(na1472_1), .IN1(1'b1), .IN2(~na399_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na417_2), .IN8(na416_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x45y103     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1475_1 ( .OUT(na1475_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na419_1), .IN8(na418_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x44y113     80'h00_0018_00_0000_0888_1533
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1476_1 ( .OUT(na1476_1), .IN1(1'b1), .IN2(~na1136_1), .IN3(1'b1), .IN4(~na1143_1), .IN5(~na1141_1), .IN6(1'b1), .IN7(~na1133_1),
                      .IN8(~na1138_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x46y109     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1478_4 ( .OUT(na1478_2), .IN1(na265_1), .IN2(1'b1), .IN3(na14_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y110     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1479_1 ( .OUT(na1479_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na422_1), .IN8(na421_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y116     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1480_1 ( .OUT(na1480_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1136_1), .IN7(na1701_2), .IN8(na1481_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x44y116     80'h00_0018_00_0040_0C64_3500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1481_1 ( .OUT(na1481_1), .IN1(1'b0), .IN2(1'b1), .IN3(~na1133_1), .IN4(1'b0), .IN5(~na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1138_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y111     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1482_1 ( .OUT(na1482_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na425_1), .IN8(na421_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x54y116     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1483_1 ( .OUT(na1483_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na426_1), .IN7(1'b1), .IN8(na1143_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x48y116     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1484_4 ( .OUT(na1484_2), .IN1(1'b1), .IN2(~na1136_1), .IN3(na1133_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y109     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1486_1 ( .OUT(na1486_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na428_1), .IN8(na427_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y115     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1487_1 ( .OUT(na1487_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na429_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y109     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1489_1 ( .OUT(na1489_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na431_1), .IN8(na427_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y117     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1490_1 ( .OUT(na1490_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na73_1), .IN7(1'b1), .IN8(na1143_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x46y106     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1491_1 ( .OUT(na1491_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na432_1), .IN8(~na433_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x50y118     80'h00_0060_00_0000_0C08_FF44
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1492_4 ( .OUT(na1492_2), .IN1(~na1141_1), .IN2(na1136_1), .IN3(~na1246_1), .IN4(na1143_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y110     80'h00_0018_00_0040_0AC8_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1493_1 ( .OUT(na1493_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na432_2), .IN8(~na435_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y114     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1494_1 ( .OUT(na1494_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na110_1), .IN7(1'b1), .IN8(na1143_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x45y105     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1495_1 ( .OUT(na1495_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na437_1), .IN6(na436_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y113     80'h00_0018_00_0000_0C88_41FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1496_1 ( .OUT(na1496_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1141_1), .IN6(~na1136_1), .IN7(~na1246_1),
                      .IN8(na1143_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x44y110     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1497_1 ( .OUT(na1497_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na439_1), .IN6(na436_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x45y113     80'h00_0018_00_0000_0EEE_BAC5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1498_1 ( .OUT(na1498_1), .IN1(~na265_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1138_1), .IN5(na1371_1), .IN6(1'b0), .IN7(na1698_2),
                      .IN8(~na1143_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y115     80'h00_0018_00_0000_0888_2FC8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1500_1 ( .OUT(na1500_1), .IN1(na1141_1), .IN2(na1136_1), .IN3(1'b1), .IN4(na1138_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1133_1),
                      .IN8(~na1143_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y105     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1501_1 ( .OUT(na1501_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na442_1), .IN6(na441_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x48y118     80'h00_0060_00_0000_0C08_FF8A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1502_4 ( .OUT(na1502_2), .IN1(na1371_1), .IN2(1'b1), .IN3(na1698_2), .IN4(na1138_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x44y105     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1504_1 ( .OUT(na1504_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na446_1), .IN6(na581_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y113     80'h00_0018_00_0040_0A81_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1506_1 ( .OUT(na1506_1), .IN1(1'b1), .IN2(~na1136_1), .IN3(~na1133_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b0), .IN7(1'b0), .IN8(na1138_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y95     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1507_1 ( .OUT(na1507_1), .IN1(1'b1), .IN2(na384_1), .IN3(1'b0), .IN4(1'b0), .IN5(na451_1), .IN6(~na452_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y103     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1508_1 ( .OUT(na1508_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na454_2), .IN6(na453_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x48y117     80'h00_0018_00_0040_0C98_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1510_1 ( .OUT(na1510_1), .IN1(1'b1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1138_1), .IN5(1'b1), .IN6(na1136_1), .IN7(~na1133_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y104     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1511_1 ( .OUT(na1511_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na456_1), .IN6(~na457_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y102     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1514_1 ( .OUT(na1514_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na459_2), .IN6(~na460_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x44y111     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1515_1 ( .OUT(na1515_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na269_1), .IN7(1'b1), .IN8(~na1143_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y104     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1516_1 ( .OUT(na1516_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na462_1), .IN6(na461_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x52y114     80'h00_0060_00_0000_0C08_FF4C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1517_4 ( .OUT(na1517_2), .IN1(1'b1), .IN2(na1136_1), .IN3(~na1699_2), .IN4(na1481_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y103     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1518_1 ( .OUT(na1518_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na464_1), .IN6(na461_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x48y114     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1519_4 ( .OUT(na1519_2), .IN1(1'b1), .IN2(~na426_1), .IN3(1'b1), .IN4(~na1143_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y101     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1520_1 ( .OUT(na1520_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na465_1), .IN6(~na466_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x54y115     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1521_1 ( .OUT(na1521_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na429_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1143_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x48y97     80'h00_0060_00_0000_0C06_FF06
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1522_4 ( .OUT(na1522_2), .IN1(na467_1), .IN2(na267_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x52y102     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1524_1 ( .OUT(na1524_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na383_1), .IN6(1'b1), .IN7(1'b1), .IN8(na70_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x44y95     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1525_4 ( .OUT(na1525_2), .IN1(1'b1), .IN2(na1441_2), .IN3(1'b1), .IN4(na1172_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x46y94     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1526_1 ( .OUT(na1526_1), .IN1(1'b1), .IN2(~na384_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na478_1), .IN8(na477_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y94     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1527_1 ( .OUT(na1527_1), .IN1(1'b1), .IN2(~na384_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na482_1), .IN6(na481_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x51y95     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1528_1 ( .OUT(na1528_1), .IN1(1'b1), .IN2(~na384_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na486_1), .IN6(na485_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y95     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1529_1 ( .OUT(na1529_1), .IN1(1'b1), .IN2(na384_1), .IN3(1'b0), .IN4(1'b0), .IN5(na489_2), .IN6(~na490_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x52y100     80'h00_0018_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1530_1 ( .OUT(na1530_1), .IN1(1'b1), .IN2(~na384_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na495_1), .IN8(na494_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x41y97     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1531_1 ( .OUT(na1531_1), .IN1(1'b1), .IN2(~na1550_2), .IN3(1'b0), .IN4(1'b0), .IN5(na675_1), .IN6(na1639_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x48y88     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1532_1 ( .OUT(na1532_1), .IN1(1'b1), .IN2(na48_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1652_2), .IN6(na705_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x32y91     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1534_4 ( .OUT(na1534_2), .IN1(1'b1), .IN2(~na160_1), .IN3(1'b1), .IN4(na576_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x38y92     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1535_1 ( .OUT(na1535_1), .IN1(1'b1), .IN2(~na1563_2), .IN3(1'b0), .IN4(1'b0), .IN5(na577_1), .IN6(na578_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y109     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1537_1 ( .OUT(na1537_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na579_1), .IN6(~na1136_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x45y106     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1538_1 ( .OUT(na1538_1), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na580_1), .IN6(na581_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x1y95     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1539_4 ( .OUT(na1539_2), .IN1(1'b1), .IN2(na499_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1539_6 ( .RAM_O2(na1539_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1539_2), .COMP_OUT(1'b0) );
// C_///AND/      x77y128     80'h08_0060_00_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1540_4 ( .OUT(na1540_2), .IN1(1'b1), .IN2(~na545_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1540_6 ( .RAM_O2(na1540_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1540_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y75     80'h08_0060_00_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1541_4 ( .OUT(na1541_2), .IN1(~na546_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1541_6 ( .RAM_O2(na1541_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1541_2), .COMP_OUT(1'b0) );
// C_///AND/      x73y128     80'h08_0060_00_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1542_4 ( .OUT(na1542_2), .IN1(1'b1), .IN2(~na388_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1542_6 ( .RAM_O2(na1542_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1542_2), .COMP_OUT(1'b0) );
// C_///AND/      x85y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1543_4 ( .OUT(na1543_2), .IN1(1'b1), .IN2(1'b1), .IN3(na468_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1543_6 ( .RAM_O2(na1543_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1543_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y71     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1544_4 ( .OUT(na1544_2), .IN1(1'b1), .IN2(1'b1), .IN3(na368_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1544_6 ( .RAM_O2(na1544_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1544_2), .COMP_OUT(1'b0) );
// C_///AND/      x81y128     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1545_4 ( .OUT(na1545_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na494_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1545_6 ( .RAM_O2(na1545_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1545_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y73     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1546_4 ( .OUT(na1546_2), .IN1(na244_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1546_6 ( .RAM_O2(na1546_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1546_2), .COMP_OUT(1'b0) );
// C_///AND/      x75y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1547_4 ( .OUT(na1547_2), .IN1(1'b1), .IN2(1'b1), .IN3(na396_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1547_6 ( .RAM_O2(na1547_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1547_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y69     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1548_4 ( .OUT(na1548_2), .IN1(na218_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1548_6 ( .RAM_O2(na1548_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1548_2), .COMP_OUT(1'b0) );
// C_////Bridge      x36y103     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1549_5 ( .OUT(na1549_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na11_2) );
// C_////Bridge      x41y96     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1550_5 ( .OUT(na1550_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na13_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y87     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1551_5 ( .OUT(na1551_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na13_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y115     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1552_5 ( .OUT(na1552_2), .IN1(1'b0), .IN2(1'b0), .IN3(na17_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y108     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1553_5 ( .OUT(na1553_2), .IN1(1'b0), .IN2(1'b0), .IN3(na17_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y114     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1554_5 ( .OUT(na1554_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na19_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y105     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1555_5 ( .OUT(na1555_2), .IN1(na23_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y114     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1556_5 ( .OUT(na1556_2), .IN1(na23_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y101     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1557_5 ( .OUT(na1557_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na32_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y97     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1558_5 ( .OUT(na1558_2), .IN1(1'b0), .IN2(1'b0), .IN3(na44_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y102     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1559_5 ( .OUT(na1559_2), .IN1(1'b0), .IN2(1'b0), .IN3(na44_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y87     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1560_5 ( .OUT(na1560_2), .IN1(1'b0), .IN2(na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y90     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1561_5 ( .OUT(na1561_2), .IN1(1'b0), .IN2(na57_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y107     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1562_5 ( .OUT(na1562_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na70_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y92     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1563_5 ( .OUT(na1563_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na96_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y83     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1564_5 ( .OUT(na1564_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na138_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y84     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1565_5 ( .OUT(na1565_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na138_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y88     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1566_5 ( .OUT(na1566_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na138_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y86     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1567_5 ( .OUT(na1567_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na139_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y87     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1568_5 ( .OUT(na1568_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na139_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y94     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1569_5 ( .OUT(na1569_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na139_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x30y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1570_5 ( .OUT(na1570_2), .IN1(1'b0), .IN2(1'b0), .IN3(na141_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y85     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1571_5 ( .OUT(na1571_2), .IN1(1'b0), .IN2(1'b0), .IN3(na142_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1572_5 ( .OUT(na1572_2), .IN1(1'b0), .IN2(1'b0), .IN3(na142_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1573_5 ( .OUT(na1573_2), .IN1(1'b0), .IN2(1'b0), .IN3(na142_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y83     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1574_5 ( .OUT(na1574_2), .IN1(1'b0), .IN2(na144_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y92     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1575_5 ( .OUT(na1575_2), .IN1(1'b0), .IN2(1'b0), .IN3(na146_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y89     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1576_5 ( .OUT(na1576_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na147_2), .IN8(1'b0) );
// C_////Bridge      x31y86     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1577_5 ( .OUT(na1577_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na149_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y96     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1578_5 ( .OUT(na1578_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na155_1) );
// C_////Bridge      x34y88     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1579_5 ( .OUT(na1579_2), .IN1(1'b0), .IN2(na160_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x30y89     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1580_5 ( .OUT(na1580_2), .IN1(1'b0), .IN2(na160_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y90     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1581_5 ( .OUT(na1581_2), .IN1(1'b0), .IN2(na160_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y101     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1582_5 ( .OUT(na1582_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na164_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x30y91     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1583_5 ( .OUT(na1583_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na166_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y96     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1584_5 ( .OUT(na1584_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na167_1), .IN8(1'b0) );
// C_////Bridge      x29y93     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1585_5 ( .OUT(na1585_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na167_2), .IN8(1'b0) );
// C_////Bridge      x37y118     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1586_5 ( .OUT(na1586_2), .IN1(1'b0), .IN2(1'b0), .IN3(na176_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y120     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1587_5 ( .OUT(na1587_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na177_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y115     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1588_5 ( .OUT(na1588_2), .IN1(1'b0), .IN2(1'b0), .IN3(na180_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y113     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1589_5 ( .OUT(na1589_2), .IN1(1'b0), .IN2(na181_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y113     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1590_5 ( .OUT(na1590_2), .IN1(1'b0), .IN2(na181_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y114     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1591_5 ( .OUT(na1591_2), .IN1(na182_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y108     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1592_5 ( .OUT(na1592_2), .IN1(1'b0), .IN2(na184_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y114     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1593_5 ( .OUT(na1593_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na187_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y114     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1594_5 ( .OUT(na1594_2), .IN1(1'b0), .IN2(1'b0), .IN3(na188_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y111     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1595_5 ( .OUT(na1595_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na189_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x30y115     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1596_5 ( .OUT(na1596_2), .IN1(na192_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y115     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1597_5 ( .OUT(na1597_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na193_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y113     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1598_5 ( .OUT(na1598_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na193_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y114     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1599_5 ( .OUT(na1599_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na193_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y116     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1600_5 ( .OUT(na1600_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na193_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y114     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1601_5 ( .OUT(na1601_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na196_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y113     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1602_5 ( .OUT(na1602_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na201_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y117     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1603_5 ( .OUT(na1603_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na202_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y107     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1604_5 ( .OUT(na1604_2), .IN1(na211_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y119     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1605_5 ( .OUT(na1605_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na215_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y115     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1606_5 ( .OUT(na1606_2), .IN1(na217_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y96     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1607_5 ( .OUT(na1607_2), .IN1(1'b0), .IN2(na219_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y100     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1608_5 ( .OUT(na1608_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na219_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x30y104     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1609_5 ( .OUT(na1609_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na231_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y110     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1610_5 ( .OUT(na1610_2), .IN1(1'b0), .IN2(na233_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y109     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1611_5 ( .OUT(na1611_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na234_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y107     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1612_5 ( .OUT(na1612_2), .IN1(1'b0), .IN2(1'b0), .IN3(na241_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y100     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1613_5 ( .OUT(na1613_2), .IN1(1'b0), .IN2(1'b0), .IN3(na250_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y103     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1614_5 ( .OUT(na1614_2), .IN1(1'b0), .IN2(1'b0), .IN3(na251_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y94     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1615_5 ( .OUT(na1615_2), .IN1(1'b0), .IN2(na256_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y114     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1616_5 ( .OUT(na1616_2), .IN1(na265_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y91     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1617_5 ( .OUT(na1617_2), .IN1(1'b0), .IN2(1'b0), .IN3(na276_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y106     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1618_5 ( .OUT(na1618_2), .IN1(1'b0), .IN2(1'b0), .IN3(na276_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y101     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1619_5 ( .OUT(na1619_2), .IN1(1'b0), .IN2(na288_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y113     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1620_5 ( .OUT(na1620_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na291_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y106     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1621_5 ( .OUT(na1621_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na292_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y99     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1622_5 ( .OUT(na1622_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na292_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y111     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1623_5 ( .OUT(na1623_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na293_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y116     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1624_5 ( .OUT(na1624_2), .IN1(na297_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y118     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1625_5 ( .OUT(na1625_2), .IN1(na297_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y111     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1626_5 ( .OUT(na1626_2), .IN1(1'b0), .IN2(1'b0), .IN3(na298_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y115     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1627_5 ( .OUT(na1627_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na299_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y113     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1628_5 ( .OUT(na1628_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na300_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y113     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1629_5 ( .OUT(na1629_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na300_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y85     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1630_5 ( .OUT(na1630_2), .IN1(na311_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y96     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1631_5 ( .OUT(na1631_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na323_1) );
// C_////Bridge      x51y96     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1632_5 ( .OUT(na1632_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na331_1), .IN8(1'b0) );
// C_////Bridge      x44y87     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1633_5 ( .OUT(na1633_2), .IN1(1'b0), .IN2(na337_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y86     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1634_5 ( .OUT(na1634_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na343_1) );
// C_////Bridge      x47y86     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1635_5 ( .OUT(na1635_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na343_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y99     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1636_5 ( .OUT(na1636_2), .IN1(1'b0), .IN2(na366_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y96     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1637_5 ( .OUT(na1637_2), .IN1(1'b0), .IN2(na366_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y96     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1638_5 ( .OUT(na1638_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na367_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y96     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1639_5 ( .OUT(na1639_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na367_2) );
// C_////Bridge      x32y104     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1640_5 ( .OUT(na1640_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na371_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y95     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1641_5 ( .OUT(na1641_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na383_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y92     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1642_5 ( .OUT(na1642_2), .IN1(1'b0), .IN2(na399_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y90     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1643_5 ( .OUT(na1643_2), .IN1(na412_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y90     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1644_5 ( .OUT(na1644_2), .IN1(na412_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y94     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1645_5 ( .OUT(na1645_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na416_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y92     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1646_5 ( .OUT(na1646_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na420_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y97     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1647_5 ( .OUT(na1647_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na420_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y89     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1648_5 ( .OUT(na1648_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na448_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y88     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1649_5 ( .OUT(na1649_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na467_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y99     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1650_5 ( .OUT(na1650_2), .IN1(1'b0), .IN2(na470_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y107     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1651_5 ( .OUT(na1651_2), .IN1(1'b0), .IN2(na470_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y87     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1652_5 ( .OUT(na1652_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na497_2), .IN8(1'b0) );
// C_////Bridge      x35y109     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1653_5 ( .OUT(na1653_2), .IN1(1'b0), .IN2(1'b0), .IN3(na498_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y110     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1654_5 ( .OUT(na1654_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na535_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y113     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1655_5 ( .OUT(na1655_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na679_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y109     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1656_5 ( .OUT(na1656_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na681_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y107     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1657_5 ( .OUT(na1657_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na681_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y117     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1658_5 ( .OUT(na1658_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na683_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y95     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1659_5 ( .OUT(na1659_2), .IN1(na685_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y98     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1660_5 ( .OUT(na1660_2), .IN1(na685_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y95     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1661_5 ( .OUT(na1661_2), .IN1(na685_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y100     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1662_5 ( .OUT(na1662_2), .IN1(na685_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y102     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1663_5 ( .OUT(na1663_2), .IN1(1'b0), .IN2(na687_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y100     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1664_5 ( .OUT(na1664_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na687_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y103     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1665_5 ( .OUT(na1665_2), .IN1(na689_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y98     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1666_5 ( .OUT(na1666_2), .IN1(na689_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y112     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1667_5 ( .OUT(na1667_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na711_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y114     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1668_5 ( .OUT(na1668_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na713_1), .IN8(1'b0) );
// C_////Bridge      x51y104     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1669_5 ( .OUT(na1669_2), .IN1(1'b0), .IN2(1'b0), .IN3(na713_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y112     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1670_5 ( .OUT(na1670_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na715_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y110     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1671_5 ( .OUT(na1671_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na728_1) );
// C_////Bridge      x27y117     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1672_5 ( .OUT(na1672_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na750_1) );
// C_////Bridge      x25y117     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1673_5 ( .OUT(na1673_2), .IN1(1'b0), .IN2(1'b0), .IN3(na752_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y111     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1674_5 ( .OUT(na1674_2), .IN1(1'b0), .IN2(1'b0), .IN3(na755_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y105     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1675_5 ( .OUT(na1675_2), .IN1(na774_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y109     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1676_5 ( .OUT(na1676_2), .IN1(na774_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y111     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1677_5 ( .OUT(na1677_2), .IN1(1'b0), .IN2(na776_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y112     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1678_5 ( .OUT(na1678_2), .IN1(1'b0), .IN2(na776_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y109     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1679_5 ( .OUT(na1679_2), .IN1(1'b0), .IN2(na776_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x30y112     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1680_5 ( .OUT(na1680_2), .IN1(1'b0), .IN2(na776_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y109     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1681_5 ( .OUT(na1681_2), .IN1(na778_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y101     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1682_5 ( .OUT(na1682_2), .IN1(na785_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y114     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1683_5 ( .OUT(na1683_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na796_1), .IN8(1'b0) );
// C_////Bridge      x34y116     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1684_5 ( .OUT(na1684_2), .IN1(1'b0), .IN2(1'b0), .IN3(na796_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y108     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1685_5 ( .OUT(na1685_2), .IN1(1'b0), .IN2(1'b0), .IN3(na800_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y93     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1686_5 ( .OUT(na1686_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na803_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y89     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1687_5 ( .OUT(na1687_2), .IN1(1'b0), .IN2(1'b0), .IN3(na805_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y87     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1688_5 ( .OUT(na1688_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na805_2), .IN8(1'b0) );
// C_////Bridge      x37y91     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1689_5 ( .OUT(na1689_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na807_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y93     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1690_5 ( .OUT(na1690_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na811_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y93     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1691_5 ( .OUT(na1691_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na820_1) );
// C_////Bridge      x31y115     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1692_5 ( .OUT(na1692_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na842_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y117     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1693_5 ( .OUT(na1693_2), .IN1(1'b0), .IN2(1'b0), .IN3(na844_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y113     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1694_5 ( .OUT(na1694_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na920_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y117     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1695_5 ( .OUT(na1695_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1030_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y106     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1696_5 ( .OUT(na1696_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1133_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y117     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1697_5 ( .OUT(na1697_2), .IN1(1'b0), .IN2(na1136_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y113     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1698_5 ( .OUT(na1698_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1141_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y113     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1699_5 ( .OUT(na1699_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1143_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y114     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1700_5 ( .OUT(na1700_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1143_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1701_5 ( .OUT(na1701_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1143_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y103     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1702_5 ( .OUT(na1702_2), .IN1(1'b0), .IN2(na1194_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y92     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1703_5 ( .OUT(na1703_2), .IN1(na1228_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y115     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1704_5 ( .OUT(na1704_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1274_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y87     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1705_5 ( .OUT(na1705_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1301_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y97     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1706_5 ( .OUT(na1706_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1359_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y102     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1707_5 ( .OUT(na1707_2), .IN1(na1363_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x30y98     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1708_5 ( .OUT(na1708_2), .IN1(na1363_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
endmodule
