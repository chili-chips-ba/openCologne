mem['h0000] = 32'h00001517;
mem['h0001] = 32'hC1C50513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'hFF060613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFD050513;
mem['h000E] = 32'h84818593;
mem['h000F] = 32'h00B55863;
mem['h0010] = 32'h00052023;
mem['h0011] = 32'h00450513;
mem['h0012] = 32'hFEB54CE3;
mem['h0013] = 32'h10008117;
mem['h0014] = 32'hFB410113;
mem['h0015] = 32'h10000197;
mem['h0016] = 32'h7AC18193;
mem['h0017] = 32'h00A54533;
mem['h0018] = 32'h00B5C5B3;
mem['h0019] = 32'h00C64633;
mem['h001A] = 32'h248000EF;
mem['h001B] = 32'h0000006F;
mem['h001C] = 32'hFD010113;
mem['h001D] = 32'h02812623;
mem['h001E] = 32'h03010413;
mem['h001F] = 32'hFCA42E23;
mem['h0020] = 32'hFCB42C23;
mem['h0021] = 32'hFCC42A23;
mem['h0022] = 32'hFE042623;
mem['h0023] = 32'h0300006F;
mem['h0024] = 32'hFD842703;
mem['h0025] = 32'hFEC42783;
mem['h0026] = 32'h00F70733;
mem['h0027] = 32'hFDC42683;
mem['h0028] = 32'hFEC42783;
mem['h0029] = 32'h00F687B3;
mem['h002A] = 32'h00074703;
mem['h002B] = 32'h00E78023;
mem['h002C] = 32'hFEC42783;
mem['h002D] = 32'h00178793;
mem['h002E] = 32'hFEF42623;
mem['h002F] = 32'hFEC42703;
mem['h0030] = 32'hFD442783;
mem['h0031] = 32'hFCF766E3;
mem['h0032] = 32'h00000013;
mem['h0033] = 32'h00078513;
mem['h0034] = 32'h02C12403;
mem['h0035] = 32'h03010113;
mem['h0036] = 32'h00008067;
mem['h0037] = 32'hFE010113;
mem['h0038] = 32'h00812E23;
mem['h0039] = 32'h02010413;
mem['h003A] = 32'hFEA42623;
mem['h003B] = 32'hFEB42423;
mem['h003C] = 32'h01C0006F;
mem['h003D] = 32'hFEC42783;
mem['h003E] = 32'h00178793;
mem['h003F] = 32'hFEF42623;
mem['h0040] = 32'hFE842783;
mem['h0041] = 32'h00178793;
mem['h0042] = 32'hFEF42423;
mem['h0043] = 32'hFEC42783;
mem['h0044] = 32'h0007C703;
mem['h0045] = 32'hFE842783;
mem['h0046] = 32'h0007C783;
mem['h0047] = 32'h00F71863;
mem['h0048] = 32'hFEC42783;
mem['h0049] = 32'h0007C783;
mem['h004A] = 32'hFC0796E3;
mem['h004B] = 32'hFEC42783;
mem['h004C] = 32'h0007C783;
mem['h004D] = 32'h00078713;
mem['h004E] = 32'hFE842783;
mem['h004F] = 32'h0007C783;
mem['h0050] = 32'h40F707B3;
mem['h0051] = 32'h00078513;
mem['h0052] = 32'h01C12403;
mem['h0053] = 32'h02010113;
mem['h0054] = 32'h00008067;
mem['h0055] = 32'hFD010113;
mem['h0056] = 32'h02812623;
mem['h0057] = 32'h03010413;
mem['h0058] = 32'hFCA42E23;
mem['h0059] = 32'hFDC42783;
mem['h005A] = 32'h00279793;
mem['h005B] = 32'hFEF42623;
mem['h005C] = 32'hFEC42703;
mem['h005D] = 32'hFDC42783;
mem['h005E] = 32'h40F707B3;
mem['h005F] = 32'hFEF42623;
mem['h0060] = 32'hFEC42783;
mem['h0061] = 32'h00078513;
mem['h0062] = 32'h02C12403;
mem['h0063] = 32'h03010113;
mem['h0064] = 32'h00008067;
mem['h0065] = 32'hFE010113;
mem['h0066] = 32'h00812E23;
mem['h0067] = 32'h02010413;
mem['h0068] = 32'h00050793;
mem['h0069] = 32'hFEF407A3;
mem['h006A] = 32'h00000013;
mem['h006B] = 32'h200007B7;
mem['h006C] = 32'h0007A783;
mem['h006D] = 32'h01F7D793;
mem['h006E] = 32'h0FF7F793;
mem['h006F] = 32'hFE0798E3;
mem['h0070] = 32'h200007B7;
mem['h0071] = 32'hFEF44703;
mem['h0072] = 32'h00E78023;
mem['h0073] = 32'h00000013;
mem['h0074] = 32'h01C12403;
mem['h0075] = 32'h02010113;
mem['h0076] = 32'h00008067;
mem['h0077] = 32'hFD010113;
mem['h0078] = 32'h02112623;
mem['h0079] = 32'h02812423;
mem['h007A] = 32'h03010413;
mem['h007B] = 32'hFCA42E23;
mem['h007C] = 32'hFCB42C23;
mem['h007D] = 32'hFD842783;
mem['h007E] = 32'hFFF78793;
mem['h007F] = 32'h00279793;
mem['h0080] = 32'hFEF42623;
mem['h0081] = 32'h0380006F;
mem['h0082] = 32'hFEC42783;
mem['h0083] = 32'hFDC42703;
mem['h0084] = 32'h00F757B3;
mem['h0085] = 32'h00F7F793;
mem['h0086] = 32'h00001737;
mem['h0087] = 32'hBD870713;
mem['h0088] = 32'h00F707B3;
mem['h0089] = 32'h0007C783;
mem['h008A] = 32'h00078513;
mem['h008B] = 32'hF69FF0EF;
mem['h008C] = 32'hFEC42783;
mem['h008D] = 32'hFFC78793;
mem['h008E] = 32'hFEF42623;
mem['h008F] = 32'hFEC42783;
mem['h0090] = 32'hFC07D4E3;
mem['h0091] = 32'h00000013;
mem['h0092] = 32'h00000013;
mem['h0093] = 32'h02C12083;
mem['h0094] = 32'h02812403;
mem['h0095] = 32'h03010113;
mem['h0096] = 32'h00008067;
mem['h0097] = 32'hFE010113;
mem['h0098] = 32'h00112E23;
mem['h0099] = 32'h00812C23;
mem['h009A] = 32'h02010413;
mem['h009B] = 32'hFEA42623;
mem['h009C] = 32'h01C0006F;
mem['h009D] = 32'hFEC42783;
mem['h009E] = 32'h00178713;
mem['h009F] = 32'hFEE42623;
mem['h00A0] = 32'h0007C783;
mem['h00A1] = 32'h00078513;
mem['h00A2] = 32'hF0DFF0EF;
mem['h00A3] = 32'hFEC42783;
mem['h00A4] = 32'h0007C783;
mem['h00A5] = 32'hFE0790E3;
mem['h00A6] = 32'h00000013;
mem['h00A7] = 32'h00000013;
mem['h00A8] = 32'h01C12083;
mem['h00A9] = 32'h01812403;
mem['h00AA] = 32'h02010113;
mem['h00AB] = 32'h00008067;
mem['h00AC] = 32'hFE010113;
mem['h00AD] = 32'h00112E23;
mem['h00AE] = 32'h00812C23;
mem['h00AF] = 32'h02010413;
mem['h00B0] = 32'h200007B7;
mem['h00B1] = 32'h00300713;
mem['h00B2] = 32'h00E78C23;
mem['h00B3] = 32'h200007B7;
mem['h00B4] = 32'h0047A783;
mem['h00B5] = 32'h00078F13;
mem['h00B6] = 32'h000F0713;
mem['h00B7] = 32'h800007B7;
mem['h00B8] = 32'h00F777B3;
mem['h00B9] = 32'h28078863;
mem['h00BA] = 32'h000F0713;
mem['h00BB] = 32'h400007B7;
mem['h00BC] = 32'h00F777B3;
mem['h00BD] = 32'h00078C63;
mem['h00BE] = 32'h82018023;
mem['h00BF] = 32'h200007B7;
mem['h00C0] = 32'h00100713;
mem['h00C1] = 32'h02E78423;
mem['h00C2] = 32'h2780006F;
mem['h00C3] = 32'h0FFF7713;
mem['h00C4] = 32'h02400793;
mem['h00C5] = 32'h08F71863;
mem['h00C6] = 32'h82018793;
mem['h00C7] = 32'h0017C703;
mem['h00C8] = 32'h0FF00793;
mem['h00C9] = 32'h00F71A63;
mem['h00CA] = 32'h200007B7;
mem['h00CB] = 32'h00200713;
mem['h00CC] = 32'h02E78423;
mem['h00CD] = 32'h24C0006F;
mem['h00CE] = 32'h8201C703;
mem['h00CF] = 32'h0FF00793;
mem['h00D0] = 32'h00F71863;
mem['h00D1] = 32'h200007B7;
mem['h00D2] = 32'h00300713;
mem['h00D3] = 32'h02E78423;
mem['h00D4] = 32'hFFF00713;
mem['h00D5] = 32'h82E18023;
mem['h00D6] = 32'h80018C23;
mem['h00D7] = 32'h100007B7;
mem['h00D8] = 32'h00078793;
mem['h00D9] = 32'h000780A3;
mem['h00DA] = 32'h100007B7;
mem['h00DB] = 32'h00078793;
mem['h00DC] = 32'h00078023;
mem['h00DD] = 32'h100007B7;
mem['h00DE] = 32'h00078793;
mem['h00DF] = 32'h0007A223;
mem['h00E0] = 32'h100007B7;
mem['h00E1] = 32'h00078793;
mem['h00E2] = 32'h0007A423;
mem['h00E3] = 32'h100007B7;
mem['h00E4] = 32'h00078793;
mem['h00E5] = 32'h0007A623;
mem['h00E6] = 32'h200007B7;
mem['h00E7] = 32'h02078423;
mem['h00E8] = 32'h1E00006F;
mem['h00E9] = 32'h8201C783;
mem['h00EA] = 32'h00079A63;
mem['h00EB] = 32'h200007B7;
mem['h00EC] = 32'h00400713;
mem['h00ED] = 32'h02E78423;
mem['h00EE] = 32'h1C80006F;
mem['h00EF] = 32'h0FFF7793;
mem['h00F0] = 32'h02C00713;
mem['h00F1] = 32'h00E78E63;
mem['h00F2] = 32'h02C00713;
mem['h00F3] = 32'h14F74463;
mem['h00F4] = 32'h00A00713;
mem['h00F5] = 32'h12E78663;
mem['h00F6] = 32'h00D00713;
mem['h00F7] = 32'h12E79C63;
mem['h00F8] = 32'h100007B7;
mem['h00F9] = 32'h00078793;
mem['h00FA] = 32'h0017C703;
mem['h00FB] = 32'h00300793;
mem['h00FC] = 32'h18E7E663;
mem['h00FD] = 32'h8001AE23;
mem['h00FE] = 32'hFE0407A3;
mem['h00FF] = 32'h0440006F;
mem['h0100] = 32'h81C1A703;
mem['h0101] = 32'h00070793;
mem['h0102] = 32'h00279793;
mem['h0103] = 32'h00E787B3;
mem['h0104] = 32'h00179793;
mem['h0105] = 32'h00078693;
mem['h0106] = 32'hFEF44783;
mem['h0107] = 32'h81018713;
mem['h0108] = 32'h00F707B3;
mem['h0109] = 32'h0007C783;
mem['h010A] = 32'h00F687B3;
mem['h010B] = 32'hFD078713;
mem['h010C] = 32'h80E1AE23;
mem['h010D] = 32'hFEF44783;
mem['h010E] = 32'h00178793;
mem['h010F] = 32'hFEF407A3;
mem['h0110] = 32'h8181C783;
mem['h0111] = 32'hFEF44703;
mem['h0112] = 32'hFAF76CE3;
mem['h0113] = 32'h100007B7;
mem['h0114] = 32'h00078793;
mem['h0115] = 32'h0017C783;
mem['h0116] = 32'h00300713;
mem['h0117] = 32'h06E78663;
mem['h0118] = 32'h00300713;
mem['h0119] = 32'h06F74A63;
mem['h011A] = 32'h00200713;
mem['h011B] = 32'h04E78463;
mem['h011C] = 32'h00200713;
mem['h011D] = 32'h06F74263;
mem['h011E] = 32'h00078863;
mem['h011F] = 32'h00100713;
mem['h0120] = 32'h02E78063;
mem['h0121] = 32'h0540006F;
mem['h0122] = 32'h81C1A783;
mem['h0123] = 32'h0FF7F713;
mem['h0124] = 32'h100007B7;
mem['h0125] = 32'h00078793;
mem['h0126] = 32'h00E78023;
mem['h0127] = 32'h03C0006F;
mem['h0128] = 32'h81C1A703;
mem['h0129] = 32'h100007B7;
mem['h012A] = 32'h00078793;
mem['h012B] = 32'h00E7A223;
mem['h012C] = 32'h0280006F;
mem['h012D] = 32'h81C1A703;
mem['h012E] = 32'h100007B7;
mem['h012F] = 32'h00078793;
mem['h0130] = 32'h00E7A423;
mem['h0131] = 32'h0140006F;
mem['h0132] = 32'h81C1A703;
mem['h0133] = 32'h100007B7;
mem['h0134] = 32'h00078793;
mem['h0135] = 32'h00E7A623;
mem['h0136] = 32'h80018C23;
mem['h0137] = 32'h100007B7;
mem['h0138] = 32'h00078793;
mem['h0139] = 32'h0017C783;
mem['h013A] = 32'h00178793;
mem['h013B] = 32'h0FF7F713;
mem['h013C] = 32'h100007B7;
mem['h013D] = 32'h00078793;
mem['h013E] = 32'h00E780A3;
mem['h013F] = 32'h0800006F;
mem['h0140] = 32'h82018023;
mem['h0141] = 32'h82018793;
mem['h0142] = 32'hFFF00713;
mem['h0143] = 32'h00E780A3;
mem['h0144] = 32'h0700006F;
mem['h0145] = 32'h0FFF7713;
mem['h0146] = 32'h02F00793;
mem['h0147] = 32'h00E7FE63;
mem['h0148] = 32'h0FFF7713;
mem['h0149] = 32'h03900793;
mem['h014A] = 32'h00E7E863;
mem['h014B] = 32'h8181C703;
mem['h014C] = 32'h00700793;
mem['h014D] = 32'h00E7FC63;
mem['h014E] = 32'h82018023;
mem['h014F] = 32'h200007B7;
mem['h0150] = 32'h00500713;
mem['h0151] = 32'h02E78423;
mem['h0152] = 32'h0380006F;
mem['h0153] = 32'h8181C783;
mem['h0154] = 32'h00178713;
mem['h0155] = 32'h0FF77693;
mem['h0156] = 32'h80D18C23;
mem['h0157] = 32'h00078693;
mem['h0158] = 32'h0FFF7713;
mem['h0159] = 32'h81018793;
mem['h015A] = 32'h00D787B3;
mem['h015B] = 32'h00E78023;
mem['h015C] = 32'h0100006F;
mem['h015D] = 32'h00000013;
mem['h015E] = 32'h0080006F;
mem['h015F] = 32'h00000013;
mem['h0160] = 32'h82018793;
mem['h0161] = 32'h0017C783;
mem['h0162] = 32'h36078A63;
mem['h0163] = 32'h82018793;
mem['h0164] = 32'h000780A3;
mem['h0165] = 32'h100007B7;
mem['h0166] = 32'h00078793;
mem['h0167] = 32'h0017C703;
mem['h0168] = 32'h00300793;
mem['h0169] = 32'h00F70A63;
mem['h016A] = 32'h200007B7;
mem['h016B] = 32'h00600713;
mem['h016C] = 32'h02E78423;
mem['h016D] = 32'h34C0006F;
mem['h016E] = 32'h100007B7;
mem['h016F] = 32'h00078793;
mem['h0170] = 32'h0007C783;
mem['h0171] = 32'h00400713;
mem['h0172] = 32'h26E78063;
mem['h0173] = 32'h00400713;
mem['h0174] = 32'h30F74863;
mem['h0175] = 32'h00300713;
mem['h0176] = 32'h18E78C63;
mem['h0177] = 32'h00300713;
mem['h0178] = 32'h30F74063;
mem['h0179] = 32'h00100713;
mem['h017A] = 32'h00E78863;
mem['h017B] = 32'h00200713;
mem['h017C] = 32'h0CE78063;
mem['h017D] = 32'h2EC0006F;
mem['h017E] = 32'h82C1C703;
mem['h017F] = 32'h0FF00793;
mem['h0180] = 32'h00F71A63;
mem['h0181] = 32'h200007B7;
mem['h0182] = 32'h00700713;
mem['h0183] = 32'h02E78423;
mem['h0184] = 32'h2F00006F;
mem['h0185] = 32'h100007B7;
mem['h0186] = 32'h00078793;
mem['h0187] = 32'h0047A783;
mem['h0188] = 32'h00078713;
mem['h0189] = 32'h000087B7;
mem['h018A] = 32'hFFF78793;
mem['h018B] = 32'h00F777B3;
mem['h018C] = 32'h01079693;
mem['h018D] = 32'h0106D693;
mem['h018E] = 32'h00008737;
mem['h018F] = 32'hFFF70713;
mem['h0190] = 32'h00E6F733;
mem['h0191] = 32'h8241A603;
mem['h0192] = 32'hFFFF86B7;
mem['h0193] = 32'h00D676B3;
mem['h0194] = 32'h00E6E733;
mem['h0195] = 32'h82E1A223;
mem['h0196] = 32'h100007B7;
mem['h0197] = 32'h00078793;
mem['h0198] = 32'h0087A783;
mem['h0199] = 32'h0017F793;
mem['h019A] = 32'h0FF7F713;
mem['h019B] = 32'h00177713;
mem['h019C] = 32'h00F71713;
mem['h019D] = 32'h8241A603;
mem['h019E] = 32'hFFFF86B7;
mem['h019F] = 32'hFFF68693;
mem['h01A0] = 32'h00D676B3;
mem['h01A1] = 32'h00E6E733;
mem['h01A2] = 32'h82E1A223;
mem['h01A3] = 32'h200007B7;
mem['h01A4] = 32'h8241A703;
mem['h01A5] = 32'h00E7A423;
mem['h01A6] = 32'hFFF00713;
mem['h01A7] = 32'h82E18623;
mem['h01A8] = 32'h200007B7;
mem['h01A9] = 32'h00200713;
mem['h01AA] = 32'h00E78C23;
mem['h01AB] = 32'h2540006F;
mem['h01AC] = 32'h82C18793;
mem['h01AD] = 32'h0017C703;
mem['h01AE] = 32'h0FF00793;
mem['h01AF] = 32'h00F71A63;
mem['h01B0] = 32'h200007B7;
mem['h01B1] = 32'h00800713;
mem['h01B2] = 32'h02E78423;
mem['h01B3] = 32'h2340006F;
mem['h01B4] = 32'h100007B7;
mem['h01B5] = 32'h00078793;
mem['h01B6] = 32'h0047A783;
mem['h01B7] = 32'h00078713;
mem['h01B8] = 32'h000087B7;
mem['h01B9] = 32'hFFF78793;
mem['h01BA] = 32'h00F777B3;
mem['h01BB] = 32'h01079693;
mem['h01BC] = 32'h0106D693;
mem['h01BD] = 32'h00008737;
mem['h01BE] = 32'hFFF70713;
mem['h01BF] = 32'h00E6F733;
mem['h01C0] = 32'h8241A603;
mem['h01C1] = 32'hFFFF86B7;
mem['h01C2] = 32'h00D676B3;
mem['h01C3] = 32'h00E6E733;
mem['h01C4] = 32'h82E1A223;
mem['h01C5] = 32'h100007B7;
mem['h01C6] = 32'h00078793;
mem['h01C7] = 32'h0087A783;
mem['h01C8] = 32'h0017F793;
mem['h01C9] = 32'h0FF7F713;
mem['h01CA] = 32'h00177713;
mem['h01CB] = 32'h00F71713;
mem['h01CC] = 32'h8241A603;
mem['h01CD] = 32'hFFFF86B7;
mem['h01CE] = 32'hFFF68693;
mem['h01CF] = 32'h00D676B3;
mem['h01D0] = 32'h00E6E733;
mem['h01D1] = 32'h82E1A223;
mem['h01D2] = 32'h200007B7;
mem['h01D3] = 32'h8241A703;
mem['h01D4] = 32'h00E7A823;
mem['h01D5] = 32'h82C18793;
mem['h01D6] = 32'hFFF00713;
mem['h01D7] = 32'h00E780A3;
mem['h01D8] = 32'h200007B7;
mem['h01D9] = 32'h00100713;
mem['h01DA] = 32'h00E78C23;
mem['h01DB] = 32'h1940006F;
mem['h01DC] = 32'h200007B7;
mem['h01DD] = 32'h0207A783;
mem['h01DE] = 32'h01F7D793;
mem['h01DF] = 32'h0FF7F793;
mem['h01E0] = 32'h00078A63;
mem['h01E1] = 32'h200007B7;
mem['h01E2] = 32'h00900713;
mem['h01E3] = 32'h02E78423;
mem['h01E4] = 32'h1700006F;
mem['h01E5] = 32'h100007B7;
mem['h01E6] = 32'h00078793;
mem['h01E7] = 32'h0047A783;
mem['h01E8] = 32'h3FF7F793;
mem['h01E9] = 32'h01079713;
mem['h01EA] = 32'h01075713;
mem['h01EB] = 32'h3FF77713;
mem['h01EC] = 32'h01071713;
mem['h01ED] = 32'h8281A603;
mem['h01EE] = 32'hFC0106B7;
mem['h01EF] = 32'hFFF68693;
mem['h01F0] = 32'h00D676B3;
mem['h01F1] = 32'h00E6E733;
mem['h01F2] = 32'h82E1A423;
mem['h01F3] = 32'h100007B7;
mem['h01F4] = 32'h00078793;
mem['h01F5] = 32'h0087A783;
mem['h01F6] = 32'h00078713;
mem['h01F7] = 32'h000087B7;
mem['h01F8] = 32'hFFF78793;
mem['h01F9] = 32'h00F777B3;
mem['h01FA] = 32'h01079693;
mem['h01FB] = 32'h0106D693;
mem['h01FC] = 32'h00008737;
mem['h01FD] = 32'hFFF70713;
mem['h01FE] = 32'h00E6F733;
mem['h01FF] = 32'h8281A603;
mem['h0200] = 32'hFFFF86B7;
mem['h0201] = 32'h00D676B3;
mem['h0202] = 32'h00E6E733;
mem['h0203] = 32'h82E1A423;
mem['h0204] = 32'h200007B7;
mem['h0205] = 32'h8281A703;
mem['h0206] = 32'h02E7A023;
mem['h0207] = 32'h200007B7;
mem['h0208] = 32'h00078C23;
mem['h0209] = 32'h0DC0006F;
mem['h020A] = 32'h200007B7;
mem['h020B] = 32'h0247A783;
mem['h020C] = 32'h01F7D793;
mem['h020D] = 32'h0FF7F793;
mem['h020E] = 32'h00078A63;
mem['h020F] = 32'h200007B7;
mem['h0210] = 32'h00A00713;
mem['h0211] = 32'h02E78423;
mem['h0212] = 32'h0B80006F;
mem['h0213] = 32'h100007B7;
mem['h0214] = 32'h00078793;
mem['h0215] = 32'h0047A783;
mem['h0216] = 32'h3FF7F793;
mem['h0217] = 32'h01079713;
mem['h0218] = 32'h01075713;
mem['h0219] = 32'h3FF77713;
mem['h021A] = 32'h01071713;
mem['h021B] = 32'h8281A603;
mem['h021C] = 32'hFC0106B7;
mem['h021D] = 32'hFFF68693;
mem['h021E] = 32'h00D676B3;
mem['h021F] = 32'h00E6E733;
mem['h0220] = 32'h82E1A423;
mem['h0221] = 32'h100007B7;
mem['h0222] = 32'h00078793;
mem['h0223] = 32'h0087A783;
mem['h0224] = 32'h00078713;
mem['h0225] = 32'h000087B7;
mem['h0226] = 32'hFFF78793;
mem['h0227] = 32'h00F777B3;
mem['h0228] = 32'h01079693;
mem['h0229] = 32'h0106D693;
mem['h022A] = 32'h00008737;
mem['h022B] = 32'hFFF70713;
mem['h022C] = 32'h00E6F733;
mem['h022D] = 32'h8281A603;
mem['h022E] = 32'hFFFF86B7;
mem['h022F] = 32'h00D676B3;
mem['h0230] = 32'h00E6E733;
mem['h0231] = 32'h82E1A423;
mem['h0232] = 32'h200007B7;
mem['h0233] = 32'h8281A703;
mem['h0234] = 32'h02E7A223;
mem['h0235] = 32'h200007B7;
mem['h0236] = 32'h00078C23;
mem['h0237] = 32'h0240006F;
mem['h0238] = 32'h200007B7;
mem['h0239] = 32'h00B00713;
mem['h023A] = 32'h02E78423;
mem['h023B] = 32'h200007B7;
mem['h023C] = 32'h00300713;
mem['h023D] = 32'h00E78C23;
mem['h023E] = 32'h0080006F;
mem['h023F] = 32'h00000013;
mem['h0240] = 32'h82C18793;
mem['h0241] = 32'h0027D783;
mem['h0242] = 32'h0A079463;
mem['h0243] = 32'h82C1C703;
mem['h0244] = 32'h0FF00793;
mem['h0245] = 32'h04F71463;
mem['h0246] = 32'h200007B7;
mem['h0247] = 32'h0087A783;
mem['h0248] = 32'h01F7D793;
mem['h0249] = 32'h0FF7F793;
mem['h024A] = 32'h02079A63;
mem['h024B] = 32'h200007B7;
mem['h024C] = 32'h00C7A703;
mem['h024D] = 32'h82E1A823;
mem['h024E] = 32'h00100713;
mem['h024F] = 32'h82E18A23;
mem['h0250] = 32'h40000737;
mem['h0251] = 32'h82E1AE23;
mem['h0252] = 32'h82018C23;
mem['h0253] = 32'h82C18793;
mem['h0254] = 32'hFFF00713;
mem['h0255] = 32'h00E78123;
mem['h0256] = 32'h05C0006F;
mem['h0257] = 32'h82C18793;
mem['h0258] = 32'h0017C703;
mem['h0259] = 32'h0FF00793;
mem['h025A] = 32'h04F71663;
mem['h025B] = 32'h200007B7;
mem['h025C] = 32'h0107A783;
mem['h025D] = 32'h01F7D793;
mem['h025E] = 32'h0FF7F793;
mem['h025F] = 32'h02079C63;
mem['h0260] = 32'h200007B7;
mem['h0261] = 32'h0147A703;
mem['h0262] = 32'h82E1A823;
mem['h0263] = 32'h00200713;
mem['h0264] = 32'h82E18A23;
mem['h0265] = 32'h40400737;
mem['h0266] = 32'h82E1AE23;
mem['h0267] = 32'h82018C23;
mem['h0268] = 32'h82C18793;
mem['h0269] = 32'hFFF00713;
mem['h026A] = 32'h00E781A3;
mem['h026B] = 32'h0080006F;
mem['h026C] = 32'h00000013;
mem['h026D] = 32'h200007B7;
mem['h026E] = 32'h0007A783;
mem['h026F] = 32'h01F7D793;
mem['h0270] = 32'h0FF7F793;
mem['h0271] = 32'h20079663;
mem['h0272] = 32'h82C18793;
mem['h0273] = 32'h0027D783;
mem['h0274] = 32'h20078063;
mem['h0275] = 32'h8381C783;
mem['h0276] = 32'h00B00713;
mem['h0277] = 32'h1EF76063;
mem['h0278] = 32'h00279713;
mem['h0279] = 32'h000017B7;
mem['h027A] = 32'hBEC78793;
mem['h027B] = 32'h00F707B3;
mem['h027C] = 32'h0007A783;
mem['h027D] = 32'h00078067;
mem['h027E] = 32'h200007B7;
mem['h027F] = 32'h02400713;
mem['h0280] = 32'h00E78023;
mem['h0281] = 32'h1B80006F;
mem['h0282] = 32'h8341C703;
mem['h0283] = 32'h200007B7;
mem['h0284] = 32'h03070713;
mem['h0285] = 32'h0FF77713;
mem['h0286] = 32'h00E78023;
mem['h0287] = 32'h1A00006F;
mem['h0288] = 32'h200007B7;
mem['h0289] = 32'h02C00713;
mem['h028A] = 32'h00E78023;
mem['h028B] = 32'h1900006F;
mem['h028C] = 32'h8301A703;
mem['h028D] = 32'h000207B7;
mem['h028E] = 32'hFFF78793;
mem['h028F] = 32'h00F777B3;
mem['h0290] = 32'h00078513;
mem['h0291] = 32'hF10FF0EF;
mem['h0292] = 32'h00050713;
mem['h0293] = 32'h82E1AA23;
mem['h0294] = 32'h83418793;
mem['h0295] = 32'h0027C783;
mem['h0296] = 32'h00200593;
mem['h0297] = 32'h00078513;
mem['h0298] = 32'hF7CFF0EF;
mem['h0299] = 32'h1580006F;
mem['h029A] = 32'h83418793;
mem['h029B] = 32'h0017C783;
mem['h029C] = 32'h00200593;
mem['h029D] = 32'h00078513;
mem['h029E] = 32'hF64FF0EF;
mem['h029F] = 32'h1400006F;
mem['h02A0] = 32'h8341C783;
mem['h02A1] = 32'h00200593;
mem['h02A2] = 32'h00078513;
mem['h02A3] = 32'hF50FF0EF;
mem['h02A4] = 32'h12C0006F;
mem['h02A5] = 32'h200007B7;
mem['h02A6] = 32'h02C00713;
mem['h02A7] = 32'h00E78023;
mem['h02A8] = 32'h8401A223;
mem['h02A9] = 32'h1180006F;
mem['h02AA] = 32'h83C1A783;
mem['h02AB] = 32'h0007A703;
mem['h02AC] = 32'h84E1A023;
mem['h02AD] = 32'h84018793;
mem['h02AE] = 32'h0027C783;
mem['h02AF] = 32'h00200593;
mem['h02B0] = 32'h00078513;
mem['h02B1] = 32'hF18FF0EF;
mem['h02B2] = 32'h0F40006F;
mem['h02B3] = 32'h84018793;
mem['h02B4] = 32'h0017C783;
mem['h02B5] = 32'h00200593;
mem['h02B6] = 32'h00078513;
mem['h02B7] = 32'hF00FF0EF;
mem['h02B8] = 32'h0DC0006F;
mem['h02B9] = 32'h8401C783;
mem['h02BA] = 32'h00200593;
mem['h02BB] = 32'h00078513;
mem['h02BC] = 32'hEECFF0EF;
mem['h02BD] = 32'h8441A783;
mem['h02BE] = 32'h00178713;
mem['h02BF] = 32'h84E1A223;
mem['h02C0] = 32'h83C1A783;
mem['h02C1] = 32'h00478713;
mem['h02C2] = 32'h82E1AE23;
mem['h02C3] = 32'h8301A703;
mem['h02C4] = 32'h000207B7;
mem['h02C5] = 32'hFFF78793;
mem['h02C6] = 32'h00F777B3;
mem['h02C7] = 32'h00078713;
mem['h02C8] = 32'h8441A783;
mem['h02C9] = 32'h08F70663;
mem['h02CA] = 32'h00600713;
mem['h02CB] = 32'h82E18C23;
mem['h02CC] = 32'h0800006F;
mem['h02CD] = 32'h200007B7;
mem['h02CE] = 32'h00D00713;
mem['h02CF] = 32'h00E78023;
mem['h02D0] = 32'h82C18793;
mem['h02D1] = 32'h0027C703;
mem['h02D2] = 32'h0FF00793;
mem['h02D3] = 32'h00F71463;
mem['h02D4] = 32'h82018623;
mem['h02D5] = 32'h82C18793;
mem['h02D6] = 32'h0037C703;
mem['h02D7] = 32'h0FF00793;
mem['h02D8] = 32'h04F71C63;
mem['h02D9] = 32'h82C18793;
mem['h02DA] = 32'h000780A3;
mem['h02DB] = 32'h04C0006F;
mem['h02DC] = 32'h200007B7;
mem['h02DD] = 32'h00A00713;
mem['h02DE] = 32'h00E78023;
mem['h02DF] = 32'h82C18793;
mem['h02E0] = 32'h0027C703;
mem['h02E1] = 32'h0FF00793;
mem['h02E2] = 32'h00F71663;
mem['h02E3] = 32'h82C18793;
mem['h02E4] = 32'h00078123;
mem['h02E5] = 32'h82C18793;
mem['h02E6] = 32'h0037C703;
mem['h02E7] = 32'h0FF00793;
mem['h02E8] = 32'h00F71E63;
mem['h02E9] = 32'h82C18793;
mem['h02EA] = 32'h000781A3;
mem['h02EB] = 32'h0100006F;
mem['h02EC] = 32'h00000013;
mem['h02ED] = 32'h0080006F;
mem['h02EE] = 32'h00000013;
mem['h02EF] = 32'h8381C783;
mem['h02F0] = 32'h00178793;
mem['h02F1] = 32'h0FF7F713;
mem['h02F2] = 32'h82E18C23;
mem['h02F3] = 32'hF00FF06F;
mem['h02F4] = 32'h00000013;
mem['h02F5] = 32'hEF8FF06F;
mem['h02F6] = 32'h33323130;
mem['h02F7] = 32'h37363534;
mem['h02F8] = 32'h42413938;
mem['h02F9] = 32'h46454443;
mem['h02FA] = 32'h00000000;
mem['h02FB] = 32'h000009F8;
mem['h02FC] = 32'h00000A08;
mem['h02FD] = 32'h00000A20;
mem['h02FE] = 32'h00000A30;
mem['h02FF] = 32'h00000A68;
mem['h0300] = 32'h00000A80;
mem['h0301] = 32'h00000A94;
mem['h0302] = 32'h00000AA8;
mem['h0303] = 32'h00000ACC;
mem['h0304] = 32'h00000AE4;
mem['h0305] = 32'h00000B34;
mem['h0306] = 32'h00000B70;
