//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 May 2024)
//  Compile Time: 1970-01-01 00:59:59
//  Program Run:  2024-07-11 21:21:52
//  Program Call: p_r +sp -i /home/user/FPGA/Boards/GateMate/gatemate_ila/net/ila_top_synth24-07-11_21-20-57.v -o /home/user/FPGA/Boards/GateMate/gatemate_ila/p_r_out/ila_top_24-07-11_21-20-57 -sp -cCP +uCIO -ccf /home/user/FPGA/Boards/GateMate/gatemate_ila/src/ILA_top.ccf 
//  File Type:    Verilog

// Gatecount:    726
module ila_top_24-07-11_21-20-57 (clk , i_mosi_ILA , i_sclk_ILA , i_ss_ILA ,
       led , o_miso_ILA 
       ) ;

input  clk;
input  i_mosi_ILA;
input  i_sclk_ILA;
input  i_ss_ILA;

output led;
output o_miso_ILA;



wire clk;
wire led;
wire na1_1;
wire na1_1_i;
wire na1_2;
wire na1_2_i;
wire na2_2;
wire na2_2_i;
wire na3_1;
wire na3_1_i;
wire na4_1;
wire na5_1;
wire na5_1_i;
wire na6_1;
wire na6_1_i;
wire na6_2;
wire na6_2_i;
wire na7_1;
wire na7_1_i;
wire na7_2;
wire na7_2_i;
wire na8_1;
wire na8_1_i;
wire na9_1;
wire na9_1_i;
wire na11_2;
wire na12_1;
wire na13_1;
wire na13_1_i;
wire na14_1;
wire na14_1_i;
wire na15_1;
wire na15_1_i;
wire na15_2;
wire na15_2_i;
wire na17_1;
wire na17_1_i;
wire na17_2;
wire na17_2_i;
wire na19_1;
wire na19_1_i;
wire na19_2;
wire na19_2_i;
wire na20_1;
wire na20_1_i;
wire na20_2;
wire na20_2_i;
wire na21_2;
wire na21_2_i;
wire na22_1;
wire na23_1;
wire na23_1_i;
wire na24_2;
wire na25_1;
wire na25_1_i;
wire na25_2;
wire na25_2_i;
wire na27_2;
wire na27_2_i;
wire na30_1;
wire na30_1_i;
wire na31_1;
wire na31_1_i;
wire na31_2;
wire na31_2_i;
wire na32_1;
wire na32_1_i;
wire na32_2;
wire na32_2_i;
wire na33_1;
wire na33_1_i;
wire na35_1;
wire na35_1_i;
wire na36_1;
wire na38_1;
wire na38_1_i;
wire na39_1;
wire na39_1_i;
wire na40_1;
wire na40_1_i;
wire na40_2;
wire na40_2_i;
wire na41_1;
wire na41_1_i;
wire na44_1;
wire na44_1_i;
wire na44_2;
wire na44_2_i;
wire na45_1;
wire na45_1_i;
wire na47_1;
wire na47_1_i;
wire na47_2;
wire na47_2_i;
wire na49_1;
wire na49_1_i;
wire na49_2;
wire na49_2_i;
wire na51_1;
wire na51_1_i;
wire na51_2;
wire na51_2_i;
wire na53_1;
wire na53_1_i;
wire na53_2;
wire na53_2_i;
wire na55_1;
wire na55_1_i;
wire na55_2;
wire na55_2_i;
wire na57_1;
wire na57_1_i;
wire na57_2;
wire na57_2_i;
wire na60_1;
wire na60_1_i;
wire na60_2;
wire na60_2_i;
wire na62_1;
wire na62_1_i;
wire na62_2;
wire na62_2_i;
wire na64_1;
wire na64_1_i;
wire na64_2;
wire na64_2_i;
wire na67_1;
wire na67_1_i;
wire na67_2;
wire na67_2_i;
wire na69_2;
wire na69_2_i;
wire na70_1;
wire na70_1_i;
wire na73_1;
wire na73_1_i;
wire na73_2;
wire na73_2_i;
wire na76_1;
wire na76_1_i;
wire na76_2;
wire na76_2_i;
wire na78_1;
wire na79_1;
wire na79_1_i;
wire na79_2;
wire na79_2_i;
wire na80_1;
wire na80_1_i;
wire na80_2;
wire na80_2_i;
wire na81_1;
wire na83_1;
wire na83_1_i;
wire na83_2;
wire na83_2_i;
wire na84_1;
wire na84_1_i;
wire na84_2;
wire na84_2_i;
wire na85_1;
wire na85_1_i;
wire na85_2;
wire na85_2_i;
wire na87_2;
wire na87_2_i;
wire na88_2;
wire na88_2_i;
wire na90_1;
wire na90_1_i;
wire na91_1;
wire na91_1_i;
wire na91_2;
wire na91_2_i;
wire na93_1;
wire na93_1_i;
wire na94_1;
wire na94_1_i;
wire na94_2;
wire na94_2_i;
wire na97_1;
wire na97_1_i;
wire na97_2;
wire na97_2_i;
wire na99_1;
wire na99_1_i;
wire na99_2;
wire na99_2_i;
wire na100_1;
wire na100_1_i;
wire na100_2;
wire na100_2_i;
wire na102_1;
wire na102_1_i;
wire na102_2;
wire na102_2_i;
wire na103_1;
wire na103_1_i;
wire na106_1;
wire na106_1_i;
wire na107_2;
wire na107_2_i;
wire na108_1;
wire na108_1_i;
wire na110_1;
wire na110_1_i;
wire na111_1;
wire na111_1_i;
wire na112_2;
wire na112_2_i;
wire na113_1;
wire na113_1_i;
wire na114_1;
wire na114_1_i;
wire na115_2;
wire na115_2_i;
wire na116_1;
wire na117_1;
wire na117_1_i;
wire na117_2;
wire na117_2_i;
wire na118_1;
wire na118_1_i;
wire na118_2;
wire na118_2_i;
wire na119_1;
wire na119_1_i;
wire na120_1;
wire na120_1_i;
wire na121_1;
wire na121_1_i;
wire na124_1;
wire na124_1_i;
wire na125_1;
wire na125_1_i;
wire na126_1;
wire na126_1_i;
wire na127_1;
wire na127_1_i;
wire na128_1;
wire na128_1_i;
wire na129_1;
wire na129_1_i;
wire na130_1;
wire na130_1_i;
wire na131_1;
wire na131_1_i;
wire na132_1;
wire na132_1_i;
wire na133_1;
wire na133_1_i;
wire na134_1;
wire na134_1_i;
wire na135_1;
wire na135_1_i;
wire na136_1;
wire na136_1_i;
wire na137_1;
wire na137_1_i;
wire na138_1;
wire na138_1_i;
wire na140_1;
wire na140_1_i;
wire na140_2;
wire na140_2_i;
wire na141_1;
wire na141_1_i;
wire na141_2;
wire na141_2_i;
wire na144_2;
wire na145_2;
wire na145_2_i;
wire na146_1;
wire na147_2;
wire na148_1;
wire na149_1;
wire na150_2;
wire na153_1;
wire na154_2;
wire na154_2_i;
wire na155_1;
wire na156_1;
wire na156_1_i;
wire na156_2;
wire na156_2_i;
wire na157_1;
wire na158_1;
wire na158_1_i;
wire na159_1;
wire na160_1;
wire na160_1_i;
wire na161_1;
wire na162_2;
wire na162_2_i;
wire na165_1;
wire na165_2;
wire na165_4;
wire na167_1;
wire na167_2;
wire na167_4;
wire na169_1;
wire na169_2;
wire na169_4;
wire na171_1;
wire na171_2;
wire na171_4;
wire na173_1;
wire na173_2;
wire na173_4;
wire na174_1;
wire na174_2;
wire na174_4;
wire na176_1;
wire na176_2;
wire na176_4;
wire na178_1;
wire na178_2;
wire na181_1;
wire na181_2;
wire na181_4;
wire na183_1;
wire na183_2;
wire na183_4;
wire na185_1;
wire na185_2;
wire na185_4;
wire na187_1;
wire na187_2;
wire na187_4;
wire na188_1;
wire na188_4;
wire na190_1;
wire na190_2;
wire na190_4;
wire na192_1;
wire na192_2;
wire na194_1;
wire na194_2;
wire na194_4;
wire na196_1;
wire na196_2;
wire na196_4;
wire na198_1;
wire na198_2;
wire na198_4;
wire na200_1;
wire na200_2;
wire na200_4;
wire na202_1;
wire na202_2;
wire na202_4;
wire na203_1;
wire na203_4;
wire na205_1;
wire na205_2;
wire na205_4;
wire na207_1;
wire na207_2;
wire na209_1;
wire na209_2;
wire na209_4;
wire na211_1;
wire na211_2;
wire na211_4;
wire na213_1;
wire na213_2;
wire na213_4;
wire na215_1;
wire na215_2;
wire na215_4;
wire na217_1;
wire na217_2;
wire na217_4;
wire na218_1;
wire na218_4;
wire na220_1;
wire na220_2;
wire na220_4;
wire na222_1;
wire na222_2;
wire na224_1;
wire na224_2;
wire na224_4;
wire na226_1;
wire na226_2;
wire na226_4;
wire na228_1;
wire na228_2;
wire na228_4;
wire na230_1;
wire na230_2;
wire na230_4;
wire na232_1;
wire na232_2;
wire na232_4;
wire na233_1;
wire na233_4;
wire na235_1;
wire na235_2;
wire na235_4;
wire na237_1;
wire na237_2;
wire na239_1;
wire na239_2;
wire na239_4;
wire na241_1;
wire na241_2;
wire na241_4;
wire na243_1;
wire na243_2;
wire na243_4;
wire na245_1;
wire na245_2;
wire na245_4;
wire na247_1;
wire na247_2;
wire na247_4;
wire na250_1;
wire na250_2;
wire na301_1;
wire na301_1_i;
wire na302_2;
wire na302_2_i;
wire na368_2;
wire na368_2_i;
wire na389_1;
wire na390_1;
wire na391_1;
wire na392_1;
wire na393_1;
wire na396_3;
wire na396_4;
wire na396_5;
wire na396_6;
wire na397_3;
wire na397_4;
wire na397_5;
wire na397_6;
wire na402_1;
wire na403_1;
wire na404_1;
wire na405_1;
wire na406_2;
wire na407_1;
wire na407_4;
wire na408_1;
wire na408_2;
wire na409_2;
wire na410_2;
wire na411_1;
wire na411_9;
wire na412_2;
wire na413_1;
wire na414_1;
wire na415_2;
wire na416_1;
wire na417_1;
wire na418_1;
wire na419_1;
wire na419_9;
wire na420_1;
wire na421_2;
wire na422_1;
wire na423_1;
wire na424_1;
wire na425_1;
wire na426_1;
wire na427_1;
wire na428_1;
wire na429_1;
wire na430_1;
wire na431_1;
wire na432_1;
wire na433_1;
wire na434_1;
wire na435_1;
wire na436_1;
wire na437_1;
wire na438_1;
wire na439_1;
wire na440_1;
wire na441_1;
wire na442_1;
wire na443_1;
wire na444_1;
wire na445_1;
wire na445_9;
wire na446_1;
wire na447_2;
wire na448_1;
wire na449_1;
wire na450_1;
wire na451_1;
wire na452_1;
wire na453_1;
wire na454_1;
wire na455_1;
wire na456_1;
wire na457_1;
wire na458_1;
wire na458_9;
wire na459_2;
wire na460_1;
wire na460_9;
wire na461_2;
wire na462_1;
wire na463_1;
wire na463_9;
wire na464_1;
wire na465_1;
wire na466_1;
wire na467_1;
wire na468_2;
wire na469_1;
wire na470_1;
wire na471_1;
wire na471_9;
wire na472_2;
wire na473_1;
wire na473_9;
wire na474_2;
wire na475_1;
wire na476_1;
wire na477_1;
wire na478_1;
wire na479_1;
wire na480_1;
wire na481_1;
wire na481_9;
wire na482_2;
wire na483_2;
wire na484_1;
wire na484_9;
wire na485_2;
wire na486_1;
wire na487_2;
wire na488_2;
wire na489_1;
wire na489_9;
wire na490_2;
wire na491_1;
wire na491_9;
wire na492_2;
wire na493_1;
wire na493_9;
wire na494_2;
wire na495_1;
wire na495_9;
wire na496_2;
wire na497_1;
wire na497_9;
wire na498_2;
wire na499_1;
wire na499_9;
wire na500_2;
wire na501_1;
wire na501_9;
wire na502_2;
wire na503_1;
wire na503_9;
wire na504_2;
wire na505_1;
wire na505_9;
wire na506_2;
wire na507_1;
wire na507_9;
wire na508_2;
wire na509_1;
wire na509_9;
wire na510_2;
wire na511_1;
wire na511_9;
wire na512_2;
wire na513_1;
wire na513_9;
wire na514_2;
wire na515_1;
wire na515_9;
wire na516_2;
wire na517_1;
wire na517_9;
wire na518_2;
wire na519_1;
wire na519_9;
wire na520_2;
wire na521_1;
wire na521_9;
wire na522_2;
wire na523_1;
wire na523_9;
wire na524_2;
wire na525_1;
wire na525_9;
wire na526_2;
wire na527_1;
wire na527_9;
wire na528_2;
wire na529_1;
wire na529_9;
wire na530_2;
wire na531_1;
wire na531_9;
wire na532_2;
wire na533_1;
wire na533_9;
wire na534_2;
wire na535_1;
wire na535_9;
wire na536_2;
wire na537_1;
wire na537_9;
wire na538_2;
wire na539_1;
wire na539_9;
wire na540_2;
wire na541_1;
wire na541_9;
wire na542_2;
wire na543_1;
wire na543_9;
wire na544_2;
wire na545_1;
wire na545_9;
wire na546_2;
wire na547_1;
wire na547_9;
wire na548_2;
wire na549_1;
wire na549_9;
wire na550_2;
wire na551_1;
wire na551_9;
wire na552_2;
wire na553_1;
wire na553_9;
wire na554_2;
wire na555_1;
wire na555_9;
wire na556_2;
wire na557_1;
wire na557_9;
wire na558_2;
wire na559_1;
wire na559_9;
wire na560_2;
wire na561_1;
wire na561_9;
wire na562_2;
wire na563_1;
wire na563_9;
wire na564_2;
wire na565_1;
wire na565_9;
wire na566_2;
wire na567_1;
wire na567_9;
wire na568_2;
wire na569_1;
wire na569_9;
wire na570_2;
wire na571_1;
wire na571_9;
wire na572_2;
wire na573_1;
wire na573_9;
wire na574_2;
wire na575_1;
wire na575_9;
wire na576_2;
wire na577_1;
wire na578_2;
wire na579_1;
wire na580_1;
wire na580_9;
wire na581_2;
wire na582_2;
wire na583_1;
wire na583_9;
wire na584_2;
wire na585_1;
wire na585_9;
wire na586_2;
wire na587_1;
wire na587_9;
wire na588_2;
wire na589_1;
wire na589_9;
wire na590_2;
wire na591_1;
wire na591_9;
wire na592_2;
wire na593_1;
wire na593_9;
wire na594_2;
wire na595_1;
wire na595_9;
wire na596_2;
wire na597_1;
wire na597_9;
wire na598_2;
wire na599_1;
wire na599_9;
wire na600_2;
wire na601_1;
wire na601_9;
wire na602_2;
wire na603_1;
wire na603_9;
wire na604_2;
wire na605_1;
wire na605_9;
wire na606_2;
wire na607_1;
wire na607_9;
wire na608_2;
wire na609_1;
wire na609_9;
wire na610_2;
wire na611_1;
wire na611_9;
wire na612_2;
wire na613_1;
wire na613_9;
wire na614_2;
wire na615_1;
wire na615_9;
wire na616_2;
wire na617_1;
wire na617_9;
wire na618_2;
wire na619_1;
wire na619_9;
wire na620_2;
wire na621_1;
wire na621_9;
wire na622_2;
wire na623_1;
wire na623_9;
wire na624_2;
wire na625_1;
wire na625_9;
wire na626_2;
wire na627_1;
wire na627_9;
wire na628_2;
wire na629_1;
wire na629_9;
wire na630_2;
wire na631_1;
wire na631_9;
wire na632_2;
wire na633_1;
wire na633_9;
wire na634_2;
wire na635_1;
wire na635_9;
wire na636_2;
wire na637_1;
wire na637_9;
wire na638_2;
wire na639_1;
wire na639_9;
wire na640_2;
wire na641_1;
wire na641_9;
wire na642_2;
wire na643_1;
wire na643_9;
wire na644_2;
wire na645_1;
wire na645_9;
wire na646_2;
wire na647_1;
wire na647_9;
wire na648_2;
wire na649_1;
wire na649_9;
wire na650_2;
wire na651_1;
wire na651_9;
wire na652_2;
wire na653_1;
wire na653_9;
wire na654_2;
wire na655_1;
wire na655_9;
wire na656_2;
wire na657_1;
wire na657_9;
wire na658_2;
wire na659_1;
wire na659_9;
wire na660_2;
wire na661_1;
wire na661_9;
wire na662_2;
wire na663_1;
wire na663_9;
wire na664_2;
wire na665_1;
wire na665_9;
wire na666_2;
wire na667_1;
wire na667_9;
wire na668_2;
wire na669_1;
wire na669_9;
wire na670_2;
wire na671_1;
wire na671_9;
wire na672_2;
wire na673_1;
wire na673_9;
wire na674_2;
wire na675_1;
wire na675_9;
wire na676_2;
wire na677_1;
wire na677_9;
wire na678_2;
wire na679_1;
wire na679_9;
wire na680_2;
wire na681_1;
wire na681_9;
wire na682_2;
wire na683_1;
wire na683_9;
wire na684_2;
wire na685_1;
wire na685_9;
wire na686_2;
wire na687_1;
wire na687_9;
wire na688_2;
wire na689_1;
wire na690_2;
wire na691_1;
wire na692_1;
wire na692_9;
wire na693_2;
wire na694_2;
wire na695_1;
wire na695_9;
wire na696_2;
wire na697_1;
wire na697_9;
wire na698_2;
wire na699_1;
wire na699_9;
wire na700_2;
wire na701_1;
wire na701_9;
wire na702_2;
wire na703_1;
wire na703_9;
wire na704_2;
wire na705_1;
wire na705_9;
wire na706_2;
wire na707_1;
wire na707_9;
wire na708_2;
wire na709_1;
wire na709_9;
wire na710_2;
wire na711_1;
wire na711_9;
wire na712_2;
wire na713_1;
wire na713_9;
wire na714_2;
wire na715_1;
wire na715_9;
wire na716_2;
wire na717_1;
wire na717_9;
wire na718_2;
wire na719_1;
wire na719_9;
wire na720_2;
wire na721_1;
wire na721_9;
wire na722_2;
wire na723_1;
wire na723_9;
wire na724_2;
wire na725_1;
wire na725_9;
wire na726_2;
wire na727_1;
wire na727_9;
wire na728_2;
wire na729_1;
wire na729_9;
wire na730_2;
wire na731_1;
wire na731_9;
wire na732_2;
wire na733_1;
wire na733_9;
wire na734_2;
wire na735_1;
wire na735_9;
wire na736_2;
wire na737_1;
wire na737_9;
wire na738_2;
wire na739_1;
wire na739_9;
wire na740_2;
wire na741_1;
wire na741_9;
wire na742_2;
wire na743_1;
wire na743_9;
wire na744_2;
wire na745_1;
wire na745_9;
wire na746_2;
wire na747_1;
wire na747_9;
wire na748_2;
wire na749_1;
wire na749_9;
wire na750_2;
wire na751_1;
wire na751_9;
wire na752_2;
wire na753_1;
wire na753_9;
wire na754_2;
wire na755_1;
wire na755_9;
wire na756_2;
wire na757_1;
wire na757_9;
wire na758_2;
wire na759_1;
wire na759_9;
wire na760_2;
wire na761_1;
wire na761_9;
wire na762_2;
wire na763_1;
wire na763_9;
wire na764_2;
wire na765_1;
wire na765_9;
wire na766_2;
wire na767_1;
wire na767_9;
wire na768_2;
wire na769_1;
wire na769_9;
wire na770_2;
wire na771_1;
wire na771_9;
wire na772_2;
wire na773_1;
wire na773_9;
wire na774_2;
wire na775_1;
wire na775_9;
wire na776_2;
wire na777_1;
wire na777_9;
wire na778_2;
wire na779_1;
wire na779_9;
wire na780_2;
wire na781_1;
wire na781_9;
wire na782_2;
wire na783_1;
wire na783_9;
wire na784_2;
wire na785_1;
wire na785_9;
wire na786_2;
wire na787_1;
wire na787_9;
wire na788_2;
wire na789_1;
wire na789_9;
wire na790_2;
wire na791_1;
wire na791_9;
wire na792_2;
wire na793_1;
wire na793_9;
wire na794_2;
wire na795_1;
wire na795_9;
wire na796_2;
wire na797_1;
wire na797_9;
wire na798_2;
wire na799_1;
wire na799_9;
wire na800_2;
wire na801_1;
wire na802_2;
wire na803_1;
wire na804_1;
wire na804_9;
wire na805_2;
wire na806_2;
wire na807_1;
wire na807_9;
wire na808_2;
wire na809_1;
wire na809_9;
wire na810_2;
wire na811_1;
wire na811_9;
wire na812_2;
wire na813_1;
wire na813_9;
wire na814_2;
wire na815_1;
wire na815_9;
wire na816_2;
wire na817_1;
wire na817_9;
wire na818_2;
wire na819_1;
wire na819_9;
wire na820_2;
wire na821_1;
wire na821_9;
wire na822_2;
wire na823_1;
wire na823_9;
wire na824_2;
wire na825_1;
wire na825_9;
wire na826_2;
wire na827_1;
wire na827_9;
wire na828_2;
wire na829_1;
wire na829_9;
wire na830_2;
wire na831_1;
wire na831_9;
wire na832_2;
wire na833_1;
wire na833_9;
wire na834_2;
wire na835_1;
wire na835_9;
wire na836_2;
wire na837_1;
wire na837_9;
wire na838_2;
wire na839_1;
wire na839_9;
wire na840_2;
wire na841_1;
wire na841_9;
wire na842_2;
wire na843_1;
wire na843_9;
wire na844_2;
wire na845_1;
wire na845_9;
wire na846_2;
wire na847_1;
wire na847_9;
wire na848_2;
wire na849_1;
wire na849_9;
wire na850_2;
wire na851_1;
wire na851_9;
wire na852_2;
wire na853_1;
wire na853_9;
wire na854_2;
wire na855_1;
wire na855_9;
wire na856_2;
wire na857_1;
wire na857_9;
wire na858_2;
wire na859_1;
wire na859_9;
wire na860_2;
wire na861_1;
wire na861_9;
wire na862_2;
wire na863_1;
wire na863_9;
wire na864_2;
wire na865_1;
wire na865_9;
wire na866_2;
wire na867_1;
wire na867_9;
wire na868_2;
wire na869_1;
wire na869_9;
wire na870_2;
wire na871_1;
wire na871_9;
wire na872_2;
wire na873_1;
wire na873_9;
wire na874_2;
wire na875_1;
wire na875_9;
wire na876_2;
wire na877_1;
wire na877_9;
wire na878_2;
wire na879_1;
wire na879_9;
wire na880_2;
wire na881_1;
wire na881_9;
wire na882_2;
wire na883_1;
wire na883_9;
wire na884_2;
wire na885_1;
wire na885_9;
wire na886_2;
wire na887_1;
wire na887_9;
wire na888_2;
wire na889_1;
wire na889_9;
wire na890_2;
wire na891_1;
wire na891_9;
wire na892_2;
wire na893_1;
wire na893_9;
wire na894_2;
wire na895_1;
wire na895_9;
wire na896_2;
wire na897_1;
wire na897_9;
wire na898_2;
wire na899_1;
wire na899_9;
wire na900_2;
wire na901_1;
wire na901_9;
wire na902_2;
wire na903_1;
wire na903_9;
wire na904_2;
wire na905_1;
wire na905_9;
wire na906_2;
wire na907_1;
wire na907_9;
wire na908_2;
wire na909_1;
wire na909_9;
wire na910_2;
wire na911_1;
wire na911_9;
wire na912_2;
wire na913_1;
wire na914_2;
wire na915_1;
wire na916_2;
wire na917_2;
wire na918_2;
wire na919_2;
wire na920_2;
wire na921_2;
wire na922_2;
wire na923_2;
wire na924_2;
wire na925_2;
wire na926_2;
wire na927_2;
wire na928_2;
wire na929_2;
wire na930_2;
wire na931_2;
wire na932_2;
wire na933_2;
wire na934_2;
wire na935_2;
wire na936_2;
wire na937_2;
wire na938_2;
wire na939_2;
wire na940_2;
wire na941_2;
wire na942_2;
wire na943_2;
wire na944_2;
wire na945_2;
wire na946_2;
wire na947_2;
wire na948_2;
wire na949_2;
wire na950_2;
wire na951_2;
wire na952_2;
wire na953_2;
wire na954_2;
wire na955_2;
wire na956_2;
wire na957_2;
wire na958_2;
wire na959_2;
wire i_ss_ILA;
wire na412_10;
wire na415_10;
wire na421_10;
wire na447_10;
wire na459_10;
wire na461_10;
wire na468_10;
wire na472_10;
wire na474_10;
wire na482_10;
wire na485_10;
wire na487_10;
wire na488_10;
wire na490_10;
wire na492_10;
wire na494_10;
wire na496_10;
wire na498_10;
wire na500_10;
wire na502_10;
wire na504_10;
wire na506_10;
wire na508_10;
wire na510_10;
wire na512_10;
wire na514_10;
wire na516_10;
wire na518_10;
wire na520_10;
wire na522_10;
wire na524_10;
wire na526_10;
wire na528_10;
wire na530_10;
wire na532_10;
wire na534_10;
wire na536_10;
wire na538_10;
wire na540_10;
wire na542_10;
wire na544_10;
wire na546_10;
wire na548_10;
wire na550_10;
wire na552_10;
wire na554_10;
wire na556_10;
wire na558_10;
wire na560_10;
wire na562_10;
wire na564_10;
wire na566_10;
wire na568_10;
wire na570_10;
wire na572_10;
wire na574_10;
wire na576_10;
wire na581_10;
wire na582_10;
wire na584_10;
wire na586_10;
wire na588_10;
wire na590_10;
wire na592_10;
wire na594_10;
wire na596_10;
wire na598_10;
wire na600_10;
wire na602_10;
wire na604_10;
wire na606_10;
wire na608_10;
wire na610_10;
wire na612_10;
wire na614_10;
wire na616_10;
wire na618_10;
wire na620_10;
wire na622_10;
wire na624_10;
wire na626_10;
wire na628_10;
wire na630_10;
wire na632_10;
wire na634_10;
wire na636_10;
wire na638_10;
wire na640_10;
wire na642_10;
wire na644_10;
wire na646_10;
wire na648_10;
wire na650_10;
wire na652_10;
wire na654_10;
wire na656_10;
wire na658_10;
wire na660_10;
wire na662_10;
wire na664_10;
wire na666_10;
wire na668_10;
wire na670_10;
wire na672_10;
wire na674_10;
wire na676_10;
wire na678_10;
wire na680_10;
wire na682_10;
wire na684_10;
wire na686_10;
wire na688_10;
wire na693_10;
wire na694_10;
wire na696_10;
wire na698_10;
wire na700_10;
wire na702_10;
wire na704_10;
wire na706_10;
wire na708_10;
wire na710_10;
wire na712_10;
wire na714_10;
wire na716_10;
wire na718_10;
wire na720_10;
wire na722_10;
wire na724_10;
wire na726_10;
wire na728_10;
wire na730_10;
wire na732_10;
wire na734_10;
wire na736_10;
wire na738_10;
wire na740_10;
wire na742_10;
wire na744_10;
wire na746_10;
wire na748_10;
wire na750_10;
wire na752_10;
wire na754_10;
wire na756_10;
wire na758_10;
wire na760_10;
wire na762_10;
wire na764_10;
wire na766_10;
wire na768_10;
wire na770_10;
wire na772_10;
wire na774_10;
wire na776_10;
wire na778_10;
wire na780_10;
wire na782_10;
wire na784_10;
wire na786_10;
wire na788_10;
wire na790_10;
wire na792_10;
wire na794_10;
wire na796_10;
wire na798_10;
wire na800_10;
wire na805_10;
wire na806_10;
wire na808_10;
wire na810_10;
wire na812_10;
wire na814_10;
wire na816_10;
wire na818_10;
wire na820_10;
wire na822_10;
wire na824_10;
wire na826_10;
wire na828_10;
wire na830_10;
wire na832_10;
wire na834_10;
wire na836_10;
wire na838_10;
wire na840_10;
wire na842_10;
wire na844_10;
wire na846_10;
wire na848_10;
wire na850_10;
wire na852_10;
wire na854_10;
wire na856_10;
wire na858_10;
wire na860_10;
wire na862_10;
wire na864_10;
wire na866_10;
wire na868_10;
wire na870_10;
wire na872_10;
wire na874_10;
wire na876_10;
wire na878_10;
wire na880_10;
wire na882_10;
wire na884_10;
wire na886_10;
wire na888_10;
wire na890_10;
wire na892_10;
wire na894_10;
wire na896_10;
wire na898_10;
wire na900_10;
wire na902_10;
wire na904_10;
wire na906_10;
wire na908_10;
wire na910_10;
wire na912_10;
wire na398_118;
wire na398_119;
wire na398_120;
wire na399_118;
wire na399_119;
wire na399_120;
wire na400_118;
wire na400_119;
wire na400_120;
wire na401_118;
wire na401_119;
wire na401_120;
wire i_mosi_ILA;
wire i_sclk_ILA;
wire o_miso_ILA;

// C_ORAND/D//AND/D      x39y42     80'h00_FE00_80_0000_0C88_AE2A
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1_1 ( .OUT(na1_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na917_2), .IN6(na1_1), .IN7(na27_2), .IN8(1'b0),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1_2 ( .OUT(na1_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1_4 ( .OUT(na1_2_i), .IN1(na140_2), .IN2(1'b1), .IN3(na27_2), .IN4(~na938_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1_5 ( .OUT(na1_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1_2_i) );
// C_///AND/D      x35y38     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2_4 ( .OUT(na2_2_i), .IN1(1'b1), .IN2(na250_2), .IN3(1'b1), .IN4(na13_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2_5 ( .OUT(na2_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2_2_i) );
// C_AND/D///      x41y45     80'h00_FD00_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3_1 ( .OUT(na3_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na393_1), .IN6(1'b1), .IN7(na4_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3_2 ( .OUT(na3_1), .CLK(~na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3_1_i) );
// C_AND////      x42y41     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4_1 ( .OUT(na4_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na922_2), .IN6(1'b1), .IN7(1'b1), .IN8(na7_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x33y45     80'h00_FD00_00_0040_0C05_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a5_1 ( .OUT(na5_1_i), .IN1(na5_1), .IN2(1'b0), .IN3(na31_1), .IN4(1'b0), .IN5(na393_1), .IN6(1'b1), .IN7(na4_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5_2 ( .OUT(na5_1), .CLK(~na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5_1_i) );
// C_AND/D//AND/D      x42y44     80'h00_FE00_80_0000_0C88_8FAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6_1 ( .OUT(na6_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na27_2), .IN8(na404_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6_2 ( .OUT(na6_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6_4 ( .OUT(na6_2_i), .IN1(1'b1), .IN2(na929_2), .IN3(na429_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6_5 ( .OUT(na6_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6_2_i) );
// C_AND*/D//ICOMP*/D      x40y40     80'h00_FE00_80_0000_0387_C595
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a7_1 ( .OUT(na7_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na393_1), .IN6(1'b1), .IN7(1'b1), .IN8(na7_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a7_2 ( .OUT(na7_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na7_1_i) );
C_ICOMP    #(.CPE_CFG (9'b1_1000_0000)) 
           _a7_4 ( .OUT(na7_2_i), .IN1(na393_1), .IN2(1'b0), .IN3(~na923_2), .IN4(~na7_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a7_5 ( .OUT(na7_2), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na7_2_i) );
// C_AND/D///      x33y42     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na929_2), .IN7(na405_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a8_2 ( .OUT(na8_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na8_1_i) );
// C_ORAND/D///      x36y40     80'h00_FD00_00_0000_0888_F5EA
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a9_1 ( .OUT(na9_1_i), .IN1(na406_2), .IN2(1'b0), .IN3(na4_1), .IN4(na160_1), .IN5(~na393_1), .IN6(1'b0), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a9_2 ( .OUT(na9_1), .CLK(~na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na9_1_i) );
// C_///AND/      x39y47     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a11_4 ( .OUT(na11_2), .IN1(na158_1), .IN2(na1_1), .IN3(na156_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x42y46     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na916_2), .IN5(~na25_2), .IN6(1'b0), .IN7(~na410_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x34y56     80'h00_FE00_00_0000_0888_EF5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1_i), .IN1(1'b0), .IN2(na409_2), .IN3(~na33_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na302_2), .IN8(na13_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a13_2 ( .OUT(na13_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na13_1_i) );
// C_ORAND/D///      x35y48     80'h00_FE00_00_0000_0888_FE5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a14_1 ( .OUT(na14_1_i), .IN1(1'b0), .IN2(na409_2), .IN3(~na33_1), .IN4(1'b0), .IN5(na301_1), .IN6(na14_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a14_2 ( .OUT(na14_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na14_1_i) );
// C_AND/D//AND/D      x34y43     80'h00_FE00_80_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a15_1 ( .OUT(na15_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na413_1), .IN6(1'b1), .IN7(na27_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a15_2 ( .OUT(na15_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na15_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a15_4 ( .OUT(na15_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na27_2), .IN4(na414_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a15_5 ( .OUT(na15_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na15_2_i) );
// C_AND/D//ORAND/D      x46y42     80'h00_FE00_80_0000_0C88_82AE
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a17_1 ( .OUT(na17_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na154_2), .IN6(~na1_1), .IN7(na27_2), .IN8(na17_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a17_2 ( .OUT(na17_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na17_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a17_4 ( .OUT(na17_2_i), .IN1(na19_1), .IN2(na927_2), .IN3(na27_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a17_5 ( .OUT(na17_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na17_2_i) );
// C_AND/D//AND/D      x45y43     80'h00_FE00_80_0000_0C88_85AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a19_1 ( .OUT(na19_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na19_2), .IN6(1'b1), .IN7(na27_2), .IN8(na368_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a19_2 ( .OUT(na19_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na19_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a19_4 ( .OUT(na19_2_i), .IN1(na428_1), .IN2(1'b1), .IN3(na27_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a19_5 ( .OUT(na19_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na19_2_i) );
// C_AND/D//AND/D      x33y53     80'h00_FE00_80_0000_0C88_CA85
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a20_1 ( .OUT(na20_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na20_2), .IN6(1'b1), .IN7(1'b1), .IN8(na13_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a20_2 ( .OUT(na20_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na20_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a20_4 ( .OUT(na20_2_i), .IN1(~na44_2), .IN2(1'b1), .IN3(na111_1), .IN4(na13_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a20_5 ( .OUT(na20_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na20_2_i) );
// C_///AND/D      x38y48     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a21_4 ( .OUT(na21_2_i), .IN1(na416_1), .IN2(na14_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a21_5 ( .OUT(na21_2), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na21_2_i) );
// C_AND////      x44y48     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3_1), .IN6(na114_1), .IN7(na119_1), .IN8(na115_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x33y49     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a23_1 ( .OUT(na23_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na14_1), .IN7(na417_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a23_2 ( .OUT(na23_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na23_1_i) );
// C_///AND/      x35y49     80'h00_0060_00_0000_0C08_FF82
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a24_4 ( .OUT(na24_2), .IN1(na3_1), .IN2(~na114_1), .IN3(na119_1), .IN4(na115_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x39y41     80'h00_FE00_80_0000_0C88_3AA5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a25_1 ( .OUT(na25_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na25_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na393_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a25_2 ( .OUT(na25_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na25_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a25_4 ( .OUT(na25_2_i), .IN1(~na393_1), .IN2(1'b1), .IN3(na31_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a25_5 ( .OUT(na25_2), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na25_2_i) );
// C_///ORAND/D      x46y41     80'h00_FE00_80_0000_0C08_FFEC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a27_4 ( .OUT(na27_2_i), .IN1(1'b0), .IN2(na14_1), .IN3(na27_2), .IN4(na22_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a27_5 ( .OUT(na27_2), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na27_2_i) );
// C_ORAND/D///      x34y44     80'h00_FE00_00_0000_0888_EF5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a30_1 ( .OUT(na30_1_i), .IN1(1'b0), .IN2(na14_1), .IN3(~na156_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na90_1), .IN8(na30_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a30_2 ( .OUT(na30_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na30_1_i) );
// C_AND/D//AND/D      x42y47     80'h00_FE00_80_0000_0C88_A5F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a31_1 ( .OUT(na31_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na393_1), .IN6(1'b1), .IN7(na31_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a31_2 ( .OUT(na31_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na31_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a31_4 ( .OUT(na31_2_i), .IN1(~na393_1), .IN2(na391_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a31_5 ( .OUT(na31_2), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na31_2_i) );
// C_AND/D//AND/D      x47y41     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a32_1 ( .OUT(na32_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na422_1), .IN7(na27_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a32_2 ( .OUT(na32_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na32_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a32_4 ( .OUT(na32_2_i), .IN1(1'b1), .IN2(na929_2), .IN3(na433_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a32_5 ( .OUT(na32_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na32_2_i) );
// C_AND/D///      x34y45     80'h00_FE00_00_0000_0888_A21A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_1 ( .OUT(na33_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(~na119_1), .IN4(~na108_1), .IN5(na5_1), .IN6(~na121_1), .IN7(na120_1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a33_2 ( .OUT(na33_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na33_1_i) );
// C_AND/D///      x33y39     80'h00_FD00_00_0000_0C88_25FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a35_1 ( .OUT(na35_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na393_1), .IN6(1'b1), .IN7(na4_1), .IN8(~na36_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a35_2 ( .OUT(na35_1), .CLK(~na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na35_1_i) );
// C_MX2b////      x44y46     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1), .IN1(1'b1), .IN2(na1_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na31_2), .IN8(~na423_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x45y41     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a38_1 ( .OUT(na38_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na424_1), .IN6(1'b1), .IN7(na27_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a38_2 ( .OUT(na38_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na38_1_i) );
// C_AND/D///      x43y38     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_1 ( .OUT(na39_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na27_2), .IN8(na425_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a39_2 ( .OUT(na39_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na39_1_i) );
// C_AND/D//AND/D      x44y41     80'h00_FE00_80_0000_0C88_8FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a40_1 ( .OUT(na40_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na27_2), .IN8(na426_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a40_2 ( .OUT(na40_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na40_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a40_4 ( .OUT(na40_2_i), .IN1(na435_1), .IN2(1'b1), .IN3(na27_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a40_5 ( .OUT(na40_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na40_2_i) );
// C_AND/D///      x45y39     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a41_1 ( .OUT(na41_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na929_2), .IN7(na427_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a41_2 ( .OUT(na41_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na41_1_i) );
// C_AND/D//AND/D      x35y53     80'h00_FE00_80_0000_0C88_4AFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a44_1 ( .OUT(na44_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na44_2), .IN6(1'b1), .IN7(~na111_1), .IN8(na13_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a44_2 ( .OUT(na44_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na44_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a44_4 ( .OUT(na44_2_i), .IN1(1'b1), .IN2(na106_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a44_5 ( .OUT(na44_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na44_2_i) );
// C_AND/D///      x44y50     80'h00_FE00_00_0000_0888_4A54
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1_i), .IN1(~na5_1), .IN2(na121_1), .IN3(~na119_1), .IN4(1'b1), .IN5(na3_1), .IN6(1'b1), .IN7(~na120_1),
                    .IN8(na108_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a45_2 ( .OUT(na45_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na45_1_i) );
// C_AND/D//AND/D      x40y59     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a47_1 ( .OUT(na47_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(1'b1), .IN8(na178_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a47_2 ( .OUT(na47_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na47_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a47_4 ( .OUT(na47_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(1'b1), .IN4(na178_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a47_5 ( .OUT(na47_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na47_2_i) );
// C_AND/D//AND/D      x36y60     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a49_1 ( .OUT(na49_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(na176_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a49_2 ( .OUT(na49_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na49_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a49_4 ( .OUT(na49_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(na176_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a49_5 ( .OUT(na49_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na49_2_i) );
// C_AND/D//AND/D      x35y58     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a51_1 ( .OUT(na51_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(1'b1), .IN8(na173_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a51_2 ( .OUT(na51_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na51_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a51_4 ( .OUT(na51_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(1'b1), .IN4(na173_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a51_5 ( .OUT(na51_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na51_2_i) );
// C_AND/D//AND/D      x36y58     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a53_1 ( .OUT(na53_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(na171_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a53_2 ( .OUT(na53_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na53_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a53_4 ( .OUT(na53_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(na171_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a53_5 ( .OUT(na53_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na53_2_i) );
// C_AND/D//AND/D      x34y57     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(1'b1), .IN8(na169_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a55_2 ( .OUT(na55_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na55_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a55_4 ( .OUT(na55_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(1'b1), .IN4(na169_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a55_5 ( .OUT(na55_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na55_2_i) );
// C_AND/D//AND/D      x37y58     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a57_1 ( .OUT(na57_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(na167_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a57_2 ( .OUT(na57_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na57_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a57_4 ( .OUT(na57_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(na167_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a57_5 ( .OUT(na57_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na57_2_i) );
// C_AND/D//AND/D      x33y55     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a60_1 ( .OUT(na60_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(1'b1), .IN8(na165_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a60_2 ( .OUT(na60_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na60_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a60_4 ( .OUT(na60_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(1'b1), .IN4(na165_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a60_5 ( .OUT(na60_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na60_2_i) );
// C_AND/D//AND/D      x34y55     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a62_1 ( .OUT(na62_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(na187_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a62_2 ( .OUT(na62_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na62_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a62_4 ( .OUT(na62_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(na187_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a62_5 ( .OUT(na62_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na62_2_i) );
// C_AND/D//AND/D      x41y41     80'h00_FE00_80_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a64_1 ( .OUT(na64_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na431_1), .IN6(1'b1), .IN7(na27_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a64_2 ( .OUT(na64_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na64_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a64_4 ( .OUT(na64_2_i), .IN1(1'b1), .IN2(na929_2), .IN3(na430_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a64_5 ( .OUT(na64_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na64_2_i) );
// C_AND/D//AND/D      x33y54     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_1 ( .OUT(na67_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(1'b1), .IN8(na185_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a67_2 ( .OUT(na67_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na67_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a67_4 ( .OUT(na67_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(1'b1), .IN4(na185_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a67_5 ( .OUT(na67_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na67_2_i) );
// C_///OR/D      x43y38     80'h00_FE00_80_0000_0C0E_FF5A
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a69_4 ( .OUT(na69_2_i), .IN1(na434_1), .IN2(1'b0), .IN3(~na27_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a69_5 ( .OUT(na69_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na69_2_i) );
// C_AND/D///      x37y59     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a70_1 ( .OUT(na70_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na403_1), .IN7(1'b1), .IN8(na13_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a70_2 ( .OUT(na70_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na70_1_i) );
// C_AND/D//AND/D      x43y39     80'h00_FE00_80_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a73_1 ( .OUT(na73_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na437_1), .IN6(1'b1), .IN7(na27_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a73_2 ( .OUT(na73_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na73_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a73_4 ( .OUT(na73_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na27_2), .IN4(na438_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a73_5 ( .OUT(na73_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na73_2_i) );
// C_AND/D//AND/D      x35y56     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a76_1 ( .OUT(na76_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(na183_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a76_2 ( .OUT(na76_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na76_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a76_4 ( .OUT(na76_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(na183_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a76_5 ( .OUT(na76_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na76_2_i) );
// C_OR////      x43y47     80'h00_0018_00_0000_0CEE_C500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na137_1), .IN6(1'b0), .IN7(1'b0), .IN8(na439_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x43y43     80'h00_FE00_80_0000_0C88_8FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a79_1 ( .OUT(na79_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na27_2), .IN8(na440_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a79_2 ( .OUT(na79_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na79_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a79_4 ( .OUT(na79_2_i), .IN1(na479_1), .IN2(1'b1), .IN3(na27_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a79_5 ( .OUT(na79_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na79_2_i) );
// C_AND/D//AND/D      x35y54     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(1'b1), .IN8(na181_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a80_2 ( .OUT(na80_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na80_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a80_4 ( .OUT(na80_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(1'b1), .IN4(na181_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a80_5 ( .OUT(na80_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na80_2_i) );
// C_OR////      x41y39     80'h00_0018_00_0000_0CEE_5A00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a81_1 ( .OUT(na81_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na441_1), .IN6(1'b0), .IN7(~na937_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x35y55     80'h00_FE00_80_0000_0C88_ACF4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a83_1 ( .OUT(na83_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na409_2), .IN7(na174_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a83_2 ( .OUT(na83_1), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na83_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a83_4 ( .OUT(na83_2_i), .IN1(~na83_2), .IN2(na409_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a83_5 ( .OUT(na83_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na83_2_i) );
// C_AND/D//AND/D      x35y43     80'h00_FE00_80_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a84_1 ( .OUT(na84_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na442_1), .IN6(1'b1), .IN7(na27_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a84_2 ( .OUT(na84_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na84_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a84_4 ( .OUT(na84_2_i), .IN1(1'b1), .IN2(na929_2), .IN3(na418_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a84_5 ( .OUT(na84_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na84_2_i) );
// C_AND/D//AND/D      x47y39     80'h00_FE00_80_0000_0C88_8FAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a85_1 ( .OUT(na85_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na27_2), .IN8(na443_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a85_2 ( .OUT(na85_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na85_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a85_4 ( .OUT(na85_2_i), .IN1(1'b1), .IN2(na444_1), .IN3(na27_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a85_5 ( .OUT(na85_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na85_2_i) );
// C_///ICOMP/D      x42y42     80'h00_FE00_80_0000_0C08_FFA9
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a87_4 ( .OUT(na87_2_i), .IN1(~na931_2), .IN2(~na1_1), .IN3(~na27_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a87_5 ( .OUT(na87_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na87_2_i) );
// C_///AND/D      x34y51     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a88_4 ( .OUT(na88_2_i), .IN1(1'b1), .IN2(na409_2), .IN3(na174_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a88_5 ( .OUT(na88_2), .CLK(na250_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na88_2_i) );
// C_AND/D///      x42y51     80'h00_FE00_00_0000_0888_42A5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1_i), .IN1(~na5_1), .IN2(1'b1), .IN3(na120_1), .IN4(1'b1), .IN5(na3_1), .IN6(~na121_1), .IN7(~na119_1),
                    .IN8(na108_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a90_2 ( .OUT(na90_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na90_1_i) );
// C_AND/D//AND/D      x36y41     80'h00_FE00_80_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a91_1 ( .OUT(na91_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na446_1), .IN6(1'b1), .IN7(na27_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a91_2 ( .OUT(na91_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na91_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a91_4 ( .OUT(na91_2_i), .IN1(1'b1), .IN2(na450_1), .IN3(na27_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a91_5 ( .OUT(na91_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na91_2_i) );
// C_ICOMP/D///      x46y39     80'h00_FE00_00_0000_0C88_A6FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_1 ( .OUT(na93_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na934_2), .IN6(~na926_2), .IN7(~na27_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a93_2 ( .OUT(na93_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na93_1_i) );
// C_AND/D//AND/D      x47y38     80'h00_FE00_80_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a94_1 ( .OUT(na94_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na448_1), .IN6(1'b1), .IN7(na27_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a94_2 ( .OUT(na94_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na94_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a94_4 ( .OUT(na94_2_i), .IN1(1'b1), .IN2(na478_1), .IN3(na27_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a94_5 ( .OUT(na94_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na94_2_i) );
// C_AND/D//AND/D      x35y46     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a97_1 ( .OUT(na97_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na451_1), .IN6(1'b1), .IN7(na27_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a97_2 ( .OUT(na97_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na97_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a97_4 ( .OUT(na97_2_i), .IN1(na452_1), .IN2(1'b1), .IN3(na27_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a97_5 ( .OUT(na97_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na97_2_i) );
// C_AND/D//AND/D      x35y44     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a99_1 ( .OUT(na99_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na453_1), .IN7(na27_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a99_2 ( .OUT(na99_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na99_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a99_4 ( .OUT(na99_2_i), .IN1(1'b1), .IN2(na929_2), .IN3(na475_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a99_5 ( .OUT(na99_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na99_2_i) );
// C_AND/D//AND/D      x49y41     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a100_1 ( .OUT(na100_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na929_2), .IN7(na454_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a100_2 ( .OUT(na100_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na100_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a100_4 ( .OUT(na100_2_i), .IN1(1'b1), .IN2(na449_1), .IN3(na27_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a100_5 ( .OUT(na100_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na100_2_i) );
// C_AND/D//AND/D      x35y42     80'h00_FE00_80_0000_0C88_8FAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a102_1 ( .OUT(na102_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na27_2), .IN8(na456_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a102_2 ( .OUT(na102_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na102_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a102_4 ( .OUT(na102_2_i), .IN1(1'b1), .IN2(na929_2), .IN3(na432_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a102_5 ( .OUT(na102_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na102_2_i) );
// C_ORAND/D///      x36y33     80'h00_FD00_00_0000_0888_F5E5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_1 ( .OUT(na103_1_i), .IN1(~na457_1), .IN2(1'b0), .IN3(na4_1), .IN4(na9_1), .IN5(~na393_1), .IN6(1'b0), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a103_2 ( .OUT(na103_1), .CLK(~na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na103_1_i) );
// C_AND/D///      x33y52     80'h00_FE00_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a106_1 ( .OUT(na106_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na113_1), .IN8(na389_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a106_2 ( .OUT(na106_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na106_1_i) );
// C_///AND/D      x38y49     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a107_4 ( .OUT(na107_2_i), .IN1(1'b1), .IN2(na14_1), .IN3(1'b1), .IN4(na462_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a107_5 ( .OUT(na107_2), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na107_2_i) );
// C_MX4b/D///      x34y42     80'h00_FD00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a108_1 ( .OUT(na108_1_i), .IN1(1'b1), .IN2(~na919_2), .IN3(1'b1), .IN4(~na393_1), .IN5(1'b0), .IN6(1'b0), .IN7(na928_2),
                     .IN8(na108_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a108_2 ( .OUT(na108_1), .CLK(~na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na108_1_i) );
// C_AND/D///      x36y57     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a110_1 ( .OUT(na110_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na390_1), .IN8(na13_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a110_2 ( .OUT(na110_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na110_1_i) );
// C_MX2b/D///      x38y53     80'h00_FE00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a111_1 ( .OUT(na111_1_i), .IN1(1'b1), .IN2(~na924_2), .IN3(1'b0), .IN4(1'b0), .IN5(na44_2), .IN6(na106_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a111_2 ( .OUT(na111_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na111_1_i) );
// C_///AND/D      x38y50     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a112_4 ( .OUT(na112_2_i), .IN1(1'b1), .IN2(na465_1), .IN3(na925_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a112_5 ( .OUT(na112_2), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na112_2_i) );
// C_AND/D///      x34y47     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a113_1 ( .OUT(na113_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na466_1), .IN6(na14_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a113_2 ( .OUT(na113_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na113_1_i) );
// C_MX4a/D///      x33y46     80'h00_FE00_00_0040_0C0A_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a114_1 ( .OUT(na114_1_i), .IN1(1'b0), .IN2(na114_1), .IN3(1'b0), .IN4(na467_1), .IN5(1'b1), .IN6(na14_1), .IN7(na119_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a114_2 ( .OUT(na114_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na114_1_i) );
// C_///ICOMP/D      x42y48     80'h00_FE00_80_0000_0C08_FF6C
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a115_4 ( .OUT(na115_2_i), .IN1(1'b0), .IN2(~na14_1), .IN3(~na116_1), .IN4(na115_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a115_5 ( .OUT(na115_2), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na115_2_i) );
// C_AND////      x38y49     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a116_1 ( .OUT(na116_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3_1), .IN6(na114_1), .IN7(na119_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x33y43     80'h00_FE00_80_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a117_1 ( .OUT(na117_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na469_1), .IN6(1'b1), .IN7(na27_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a117_2 ( .OUT(na117_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na117_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a117_4 ( .OUT(na117_2_i), .IN1(1'b1), .IN2(na436_1), .IN3(na27_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a117_5 ( .OUT(na117_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na117_2_i) );
// C_AND/D//AND/D      x44y39     80'h00_FE00_80_0000_0C88_ACAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a118_1 ( .OUT(na118_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na470_1), .IN7(na27_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a118_2 ( .OUT(na118_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na118_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a118_4 ( .OUT(na118_2_i), .IN1(na420_1), .IN2(1'b1), .IN3(na27_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a118_5 ( .OUT(na118_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na118_2_i) );
// C_ORAND/D///      x42y45     80'h00_FE00_00_0000_0888_EF5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a119_1 ( .OUT(na119_1_i), .IN1(1'b0), .IN2(na14_1), .IN3(~na27_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na119_1), .IN8(na45_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a119_2 ( .OUT(na119_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na119_1_i) );
// C_MX4b/D///      x44y49     80'h00_FD00_00_0040_0A50_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a120_1 ( .OUT(na120_1_i), .IN1(na393_1), .IN2(1'b1), .IN3(~na4_1), .IN4(1'b1), .IN5(na25_2), .IN6(1'b0), .IN7(na120_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a120_2 ( .OUT(na120_1), .CLK(~na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na120_1_i) );
// C_MX4b/D///      x33y44     80'h00_FD00_00_0040_0AA0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a121_1 ( .OUT(na121_1_i), .IN1(~na393_1), .IN2(1'b1), .IN3(na4_1), .IN4(1'b1), .IN5(1'b0), .IN6(na121_1), .IN7(1'b0), .IN8(na930_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a121_2 ( .OUT(na121_1), .CLK(~na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na121_1_i) );
// C_MX2b/D///      x34y40     80'h00_F600_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a124_1 ( .OUT(na124_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na15_2), .IN8(~na124_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a124_2 ( .OUT(na124_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na124_1_i) );
// C_MX2b/D///      x35y41     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a125_1 ( .OUT(na125_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na948_2), .IN8(na194_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a125_2 ( .OUT(na125_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na125_1_i) );
// C_MX2b/D///      x37y44     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a126_1 ( .OUT(na126_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na949_2), .IN8(na194_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a126_2 ( .OUT(na126_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na126_1_i) );
// C_MX2b/D///      x42y43     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a127_1 ( .OUT(na127_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na211_1), .IN8(na942_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a127_2 ( .OUT(na127_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na127_1_i) );
// C_MX2b/D///      x39y44     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na211_2), .IN8(na943_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a128_2 ( .OUT(na128_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na128_1_i) );
// C_MX2b/D///      x37y45     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a129_1 ( .OUT(na129_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na950_2), .IN8(na198_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a129_2 ( .OUT(na129_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na129_1_i) );
// C_MX2b/D///      x38y45     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a130_1 ( .OUT(na130_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na951_2), .IN8(na198_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a130_2 ( .OUT(na130_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na130_1_i) );
// C_MX2b/D///      x39y45     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a131_1 ( .OUT(na131_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na215_1), .IN8(na944_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a131_2 ( .OUT(na131_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na131_1_i) );
// C_MX2b/D///      x37y46     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a132_1 ( .OUT(na132_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na215_2), .IN8(na945_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a132_2 ( .OUT(na132_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na132_1_i) );
// C_MX2b/D///      x38y46     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a133_1 ( .OUT(na133_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na952_2), .IN8(na202_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a133_2 ( .OUT(na133_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na133_1_i) );
// C_MX2b/D///      x37y47     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a134_1 ( .OUT(na134_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na953_2), .IN8(na202_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a134_2 ( .OUT(na134_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na134_1_i) );
// C_MX2b/D///      x38y47     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a135_1 ( .OUT(na135_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na205_1), .IN8(na940_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a135_2 ( .OUT(na135_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na135_1_i) );
// C_MX2b/D///      x37y48     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a136_1 ( .OUT(na136_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na205_2), .IN8(na941_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a136_2 ( .OUT(na136_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na136_1_i) );
// C_MX2b/D///      x35y47     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a137_1 ( .OUT(na137_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na946_2), .IN8(na192_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a137_2 ( .OUT(na137_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na137_1_i) );
// C_MX2b/D///      x37y42     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na947_2), .IN8(na192_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a138_2 ( .OUT(na138_1), .CLK(na392_1), .EN(~na146_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na138_1_i) );
// C_AND/D//AND/D      x43y41     80'h00_FE00_80_0000_0C88_ACFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a140_1 ( .OUT(na140_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na476_1), .IN7(na27_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a140_2 ( .OUT(na140_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na140_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a140_4 ( .OUT(na140_2_i), .IN1(na140_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a140_5 ( .OUT(na140_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na140_2_i) );
// C_AND/D//AND/D      x49y40     80'h00_FE00_80_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a141_1 ( .OUT(na141_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na477_1), .IN6(1'b1), .IN7(na27_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a141_2 ( .OUT(na141_1), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na141_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a141_4 ( .OUT(na141_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na27_2), .IN4(na455_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a141_5 ( .OUT(na141_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na141_2_i) );
// C_///OR/      x39y39     80'h00_0060_00_0000_0C0E_FF0D
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a144_4 ( .OUT(na144_2), .IN1(~na137_1), .IN2(na480_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x30y49     80'h00_FE00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a145_4 ( .OUT(na145_2_i), .IN1(na44_1), .IN2(1'b1), .IN3(1'b1), .IN4(na13_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a145_5 ( .OUT(na145_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na145_2_i) );
// C_ORAND////      x36y43     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a146_1 ( .OUT(na146_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na939_2), .IN6(~na1_1), .IN7(~na918_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x36y36     80'h00_0060_00_0000_0C08_FFA2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a147_4 ( .OUT(na147_2), .IN1(na932_2), .IN2(~na1_1), .IN3(na91_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x38y51     80'h00_0018_00_0000_0C88_A1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a148_1 ( .OUT(na148_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na933_2), .IN6(~na1_1), .IN7(na91_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x36y38     80'h00_0018_00_0000_0C88_A1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a149_1 ( .OUT(na149_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na932_2), .IN6(~na1_1), .IN7(na91_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x33y42     80'h00_0060_00_0000_0C08_FF51
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a150_4 ( .OUT(na150_2), .IN1(~na932_2), .IN2(~na1_1), .IN3(~na91_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x41y51     80'h00_0018_00_0040_0C05_4000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a153_1 ( .OUT(na153_1), .IN1(na20_1), .IN2(1'b0), .IN3(na145_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na107_2), .IN8(na21_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x39y49     80'h00_FE00_80_0000_0C08_FFCE
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a154_4 ( .OUT(na154_2_i), .IN1(na154_2), .IN2(na483_2), .IN3(1'b0), .IN4(na13_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a154_5 ( .OUT(na154_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na154_2_i) );
// C_MX4b////      x35y52     80'h00_0018_00_0040_0ACF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a155_1 ( .OUT(na155_1), .IN1(1'b1), .IN2(na138_1), .IN3(~na937_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na578_2), .IN8(~na957_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//ORAND/D      x40y49     80'h00_FE00_80_0000_0C88_A7EC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a156_1 ( .OUT(na156_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na78_1), .IN6(~na155_1), .IN7(na156_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a156_2 ( .OUT(na156_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na156_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a156_4 ( .OUT(na156_2_i), .IN1(1'b0), .IN2(na14_1), .IN3(na156_2), .IN4(na464_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a156_5 ( .OUT(na156_2), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na156_2_i) );
// C_MX4b////      x39y54     80'h00_0018_00_0040_0ACF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a157_1 ( .OUT(na157_1), .IN1(1'b1), .IN2(na138_1), .IN3(~na937_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na954_2), .IN8(~na801_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x43y45     80'h00_FE00_00_0000_0C88_A7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a158_1 ( .OUT(na158_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na81_1), .IN6(~na157_1), .IN7(na156_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a158_2 ( .OUT(na158_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na158_1_i) );
// C_MX2b////      x46y48     80'h00_0018_00_0040_0A54_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a159_1 ( .OUT(na159_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na486_1), .IN6(1'b0), .IN7(~na31_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x44y44     80'h00_FD00_00_0000_0888_F57E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a160_1 ( .OUT(na160_1_i), .IN1(na35_1), .IN2(na919_2), .IN3(~na4_1), .IN4(~na159_1), .IN5(~na393_1), .IN6(1'b0), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a160_2 ( .OUT(na160_1), .CLK(~na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na160_1_i) );
// C_MX4b////      x33y48     80'h00_0018_00_0040_0ACF_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a161_1 ( .OUT(na161_1), .IN1(1'b1), .IN2(na138_1), .IN3(~na937_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na579_1), .IN8(~na958_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x39y46     80'h00_FE00_80_0000_0C08_FFA7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a162_4 ( .OUT(na162_2_i), .IN1(~na144_2), .IN2(~na161_1), .IN3(na156_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a162_5 ( .OUT(na162_2), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na162_2_i) );
// C_ADDF2///ADDF2/      x36y50     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a165_1 ( .OUT(na165_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na60_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na187_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a165_4 ( .OUT(na165_2), .COUTY1(na165_4), .IN1(na60_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na60_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na187_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y51     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a167_1 ( .OUT(na167_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na57_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na165_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a167_4 ( .OUT(na167_2), .COUTY1(na167_4), .IN1(1'b1), .IN2(na57_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na57_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na165_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y52     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a169_1 ( .OUT(na169_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na55_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na167_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a169_4 ( .OUT(na169_2), .COUTY1(na169_4), .IN1(1'b0), .IN2(1'b0), .IN3(na55_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na55_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na167_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y53     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a171_1 ( .OUT(na171_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na53_2),
                     .CINX(1'b0), .CINY1(na169_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a171_4 ( .OUT(na171_2), .COUTY1(na171_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na53_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na53_2), .CINX(1'b0), .CINY1(na169_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y54     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a173_1 ( .OUT(na173_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na51_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na171_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a173_4 ( .OUT(na173_2), .COUTY1(na173_4), .IN1(1'b1), .IN2(na51_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na51_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na171_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y45     80'h00_0078_00_0020_0C66_AA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a174_1 ( .OUT(na174_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na83_2), .IN6(1'b1), .IN7(na88_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na188_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a174_4 ( .OUT(na174_2), .COUTY1(na174_4), .IN1(na83_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na83_2), .IN6(1'b1), .IN7(na88_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na188_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y55     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a176_1 ( .OUT(na176_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na49_2),
                     .CINX(1'b0), .CINY1(na173_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a176_4 ( .OUT(na176_2), .COUTY1(na176_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na49_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na49_2), .CINX(1'b0), .CINY1(na173_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y56     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a178_1 ( .OUT(na178_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na47_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na176_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a178_4 ( .OUT(na178_2), .IN1(1'b0), .IN2(1'b0), .IN3(na47_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na47_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na176_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y46     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a181_1 ( .OUT(na181_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na80_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na174_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a181_4 ( .OUT(na181_2), .COUTY1(na181_4), .IN1(1'b1), .IN2(na80_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na80_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na174_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y47     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a183_1 ( .OUT(na183_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na76_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na181_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a183_4 ( .OUT(na183_2), .COUTY1(na183_4), .IN1(1'b1), .IN2(na76_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na76_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na181_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y48     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a185_1 ( .OUT(na185_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na67_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na183_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a185_4 ( .OUT(na185_2), .COUTY1(na185_4), .IN1(1'b1), .IN2(na67_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na67_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na183_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x36y49     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a187_1 ( .OUT(na187_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na62_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na185_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a187_4 ( .OUT(na187_2), .COUTY1(na187_4), .IN1(1'b0), .IN2(1'b0), .IN3(na62_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na62_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na185_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x36y44     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a188_2 ( .OUT(na188_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a188_6 ( .COUTY1(na188_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na188_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x40y47     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a190_1 ( .OUT(na190_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na135_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na202_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a190_4 ( .OUT(na190_2), .COUTY1(na190_4), .IN1(1'b1), .IN2(na136_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na135_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na202_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x40y48     80'h00_0078_00_0020_0C66_0A0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a192_1 ( .OUT(na192_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na137_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na190_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a192_4 ( .OUT(na192_2), .IN1(1'b1), .IN2(na138_1), .IN3(1'b0), .IN4(1'b0), .IN5(na137_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na190_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x40y42     80'h00_0078_00_0020_0C66_CA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a194_1 ( .OUT(na194_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na125_1), .IN6(1'b1), .IN7(1'b1), .IN8(na124_1),
                     .CINX(1'b0), .CINY1(na203_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a194_4 ( .OUT(na194_2), .COUTY1(na194_4), .IN1(1'b1), .IN2(na126_1), .IN3(1'b0), .IN4(1'b0), .IN5(na125_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na124_1), .CINX(1'b0), .CINY1(na203_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x40y43     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a196_1 ( .OUT(na196_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na127_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na194_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a196_4 ( .OUT(na196_2), .COUTY1(na196_4), .IN1(1'b1), .IN2(na128_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na127_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na194_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x40y44     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a198_1 ( .OUT(na198_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na129_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na196_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a198_4 ( .OUT(na198_2), .COUTY1(na198_4), .IN1(1'b0), .IN2(1'b0), .IN3(na130_1), .IN4(1'b1), .IN5(na129_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na196_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x40y45     80'h00_0078_00_0020_0C66_0A0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a200_1 ( .OUT(na200_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na131_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na198_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a200_4 ( .OUT(na200_2), .COUTY1(na200_4), .IN1(1'b1), .IN2(na132_1), .IN3(1'b0), .IN4(1'b0), .IN5(na131_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na198_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x40y46     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a202_1 ( .OUT(na202_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na133_1),
                     .CINX(1'b0), .CINY1(na200_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a202_4 ( .OUT(na202_2), .COUTY1(na202_4), .IN1(na134_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na133_1), .CINX(1'b0), .CINY1(na200_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x40y41     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a203_2 ( .OUT(na203_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a203_6 ( .COUTY1(na203_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na203_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x38y43     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a205_1 ( .OUT(na205_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na97_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na217_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a205_4 ( .OUT(na205_2), .COUTY1(na205_4), .IN1(1'b1), .IN2(na97_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na97_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na217_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y44     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a207_1 ( .OUT(na207_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na91_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na205_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a207_4 ( .OUT(na207_2), .IN1(1'b0), .IN2(1'b0), .IN3(na91_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na91_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na205_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y38     80'h00_0078_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a209_1 ( .OUT(na209_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na8_1), .IN7(na15_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na218_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a209_4 ( .OUT(na209_2), .COUTY1(na209_4), .IN1(1'b0), .IN2(1'b0), .IN3(na15_1), .IN4(1'b1), .IN5(1'b1), .IN6(na8_1), .IN7(na15_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na218_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y39     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a211_1 ( .OUT(na211_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na117_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na209_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a211_4 ( .OUT(na211_2), .COUTY1(na211_4), .IN1(na117_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na117_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na209_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y40     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a213_1 ( .OUT(na213_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na102_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na211_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a213_4 ( .OUT(na213_2), .COUTY1(na213_4), .IN1(1'b1), .IN2(na102_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na102_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na211_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y41     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a215_1 ( .OUT(na215_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na84_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na213_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a215_4 ( .OUT(na215_2), .COUTY1(na215_4), .IN1(na84_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na84_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na213_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y42     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a217_1 ( .OUT(na217_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na99_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na215_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a217_4 ( .OUT(na217_2), .COUTY1(na217_4), .IN1(1'b1), .IN2(na99_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na99_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na215_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x38y37     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a218_2 ( .OUT(na218_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a218_6 ( .COUTY1(na218_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na218_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x48y42     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a220_1 ( .OUT(na220_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na6_2),
                     .CINX(1'b0), .CINY1(na232_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a220_4 ( .OUT(na220_2), .COUTY1(na220_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na6_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na6_2), .CINX(1'b0), .CINY1(na232_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y43     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a222_1 ( .OUT(na222_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na79_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na220_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a222_4 ( .OUT(na222_2), .IN1(na79_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na79_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na220_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y37     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a224_1 ( .OUT(na224_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na73_2), .IN6(1'b1), .IN7(1'b1), .IN8(na87_2),
                     .CINX(1'b0), .CINY1(na233_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a224_4 ( .OUT(na224_2), .COUTY1(na224_4), .IN1(na73_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na73_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na87_2), .CINX(1'b0), .CINY1(na233_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y38     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a226_1 ( .OUT(na226_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na118_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na224_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a226_4 ( .OUT(na226_2), .COUTY1(na226_4), .IN1(1'b0), .IN2(1'b0), .IN3(na118_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na118_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na224_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y39     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a228_1 ( .OUT(na228_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na64_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na226_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a228_4 ( .OUT(na228_2), .COUTY1(na228_4), .IN1(na64_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na64_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na226_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y40     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a230_1 ( .OUT(na230_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na40_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na228_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a230_4 ( .OUT(na230_2), .COUTY1(na230_4), .IN1(1'b0), .IN2(1'b0), .IN3(na40_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na40_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na228_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x48y41     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a232_1 ( .OUT(na232_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na41_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na230_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a232_4 ( .OUT(na232_2), .COUTY1(na232_4), .IN1(na19_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na41_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na230_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x48y36     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a233_2 ( .OUT(na233_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a233_6 ( .COUTY1(na233_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na233_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x51y41     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a235_1 ( .OUT(na235_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na69_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na247_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a235_4 ( .OUT(na235_2), .COUTY1(na235_4), .IN1(1'b1), .IN2(na39_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na69_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na247_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y42     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a237_1 ( .OUT(na237_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na38_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na235_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a237_4 ( .OUT(na237_2), .IN1(na140_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na38_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na235_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y36     80'h00_0078_00_0020_0C66_AA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a239_1 ( .OUT(na239_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na85_2), .IN6(1'b1), .IN7(na93_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na407_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a239_4 ( .OUT(na239_2), .COUTY1(na239_4), .IN1(na85_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na85_2), .IN6(1'b1), .IN7(na93_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na407_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y37     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a241_1 ( .OUT(na241_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na94_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na239_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a241_4 ( .OUT(na241_2), .COUTY1(na241_4), .IN1(1'b1), .IN2(na94_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na94_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na239_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y38     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a243_1 ( .OUT(na243_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na100_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na241_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a243_4 ( .OUT(na243_2), .COUTY1(na243_4), .IN1(na100_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na100_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na241_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y39     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a245_1 ( .OUT(na245_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na141_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na243_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a245_4 ( .OUT(na245_2), .COUTY1(na245_4), .IN1(1'b1), .IN2(na141_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na141_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na243_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y40     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a247_1 ( .OUT(na247_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na32_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na245_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a247_4 ( .OUT(na247_2), .COUTY1(na247_4), .IN1(na32_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na32_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na245_4), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0014_0016)) 
           _a250 ( .GLB0(na250_1), .GLB1(na250_2), .GLB2(_d0), .GLB3(_d1), .CLK_FB0(_d2), .CLK_FB1(_d3), .CLK_FB2(_d4), .CLK_FB3(_d5),
                   .CLK0_0(na397_6), .CLK0_90(na397_5), .CLK0_180(na397_4), .CLK0_270(na397_3), .CLK0_BYP(1'b0), .CLK1_0(na396_6),
                   .CLK1_90(na396_5), .CLK1_180(na396_4), .CLK1_270(na396_3), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0),
                   .CLK2_270(1'b0), .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0),
                   .USR_GLB0(1'b0), .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0),
                   .USR_FB3(1'b0) );
// C_AND/D///      x33y47     80'h00_FE00_00_0000_0C88_F3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a301_1 ( .OUT(na301_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na14_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a301_2 ( .OUT(na301_1), .CLK(na392_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na301_1_i) );
// C_///AND/D      x34y53     80'h00_FE00_80_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a302_4 ( .OUT(na302_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na13_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a302_5 ( .OUT(na302_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na302_2_i) );
// C_///AND/D      x46y40     80'h00_FE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a368_4 ( .OUT(na368_2_i), .IN1(na19_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a368_5 ( .OUT(na368_2), .CLK(na250_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na368_2_i) );
// C_MX4b////      x34y54     80'h00_0018_00_0040_0A70_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a389_1 ( .OUT(na389_1), .IN1(na23_1), .IN2(1'b1), .IN3(1'b1), .IN4(na112_2), .IN5(na70_1), .IN6(na2_2), .IN7(na110_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a390 ( .Y(na390_1), .I(clk) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a391 ( .Y(na391_1), .I(i_mosi_ILA) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a392 ( .Y(na392_1), .I(i_sclk_ILA) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a393 ( .Y(na393_1), .I(i_ss_ILA) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a394 ( .O(led), .A(na487_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a395 ( .O(o_miso_ILA), .A(na488_10) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_0C_08_0C_20_82)) 
           _a396 ( .USR_PLL_LOCKED_STDY(_d6), .USR_PLL_LOCKED(_d7), .CLK270(na396_3), .CLK180(na396_4), .CLK90(na396_5), .CLK0(na396_6),
                   .CLK_REF_OUT(_d8), .CLK_REF(na408_2), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_EB_08_2F_08_82)) 
           _a397 ( .USR_PLL_LOCKED_STDY(_d9), .USR_PLL_LOCKED(_d10), .CLK270(na397_3), .CLK180(na397_4), .CLK90(na397_5), .CLK0(na397_6),
                   .CLK_REF_OUT(_d11), .CLK_REF(na408_1), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_01_04_05_00_60_00_0C_00_00_00_03_13_00_00_00_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a398 ( .DOA({_d12, _d13, _d14, _d15, _d16, _d17, _d18, _d19, _d20, _d21, _d22, _d23, _d24, _d25, _d26, _d27, _d28, _d29,
                  _d30, _d31, _d32, _d33, _d34, _d35, _d36, _d37, _d38, _d39, _d40, _d41, _d42, _d43, _d44, _d45, _d46, _d47, _d48,
                  _d49, _d50, _d51}),
                   .DOAX({_d52, _d53, _d54, _d55, _d56, _d57, _d58, _d59, _d60, _d61, _d62, _d63, _d64, _d65, _d66, _d67, _d68, _d69,
                  _d70, _d71, _d72, _d73, _d74, _d75, _d76, _d77, _d78, _d79, _d80, _d81, _d82, _d83, _d84, _d85, _d86, _d87, _d88,
                  _d89, _d90, _d91}),
                   .DOB({_d92, _d93, _d94, _d95, _d96, _d97, _d98, _d99, _d100, _d101, _d102, _d103, _d104, _d105, _d106, _d107, _d108,
                  _d109, _d110, _d111, _d112, _d113, _d114, _d115, _d116, _d117, _d118, _d119, _d120, _d121, _d122, _d123, _d124, _d125,
                  _d126, _d127, _d128, na398_118, na398_119, na398_120}),
                   .DOBX({_d129, _d130, _d131, _d132, _d133, _d134, _d135, _d136, _d137, _d138, _d139, _d140, _d141, _d142, _d143,
                  _d144, _d145, _d146, _d147, _d148, _d149, _d150, _d151, _d152, _d153, _d154, _d155, _d156, _d157, _d158, _d159, _d160,
                  _d161, _d162, _d163, _d164, _d165, _d166, _d167, _d168}),
                   .ECC1B_ERRA({_d169, _d170, _d171, _d172}),
                   .ECC1B_ERRB({_d173, _d174, _d175, _d176}),
                   .ECC2B_ERRA({_d177, _d178, _d179, _d180}),
                   .ECC2B_ERRB({_d181, _d182, _d183, _d184}),
                   .FORW_CAS_WRAO(_d185), .FORW_CAS_WRBO(_d186), .FORW_CAS_BMAO(_d187), .FORW_CAS_BMBO(_d188), .FORW_CAS_RDAO(_d189),
                   .FORW_CAS_RDBO(_d190), .FORW_UADDRAO({_d191, _d192, _d193, _d194, _d195, _d196, _d197, _d198, _d199, _d200, _d201,
                  _d202, _d203, _d204, _d205, _d206}),
                   .FORW_LADDRAO({_d207, _d208, _d209, _d210, _d211, _d212, _d213, _d214, _d215, _d216, _d217, _d218, _d219, _d220,
                  _d221, _d222}),
                   .FORW_UADDRBO({_d223, _d224, _d225, _d226, _d227, _d228, _d229, _d230, _d231, _d232, _d233, _d234, _d235, _d236,
                  _d237, _d238}),
                   .FORW_LADDRBO({_d239, _d240, _d241, _d242, _d243, _d244, _d245, _d246, _d247, _d248, _d249, _d250, _d251, _d252,
                  _d253, _d254}),
                   .FORW_UA0CLKO(_d255), .FORW_UA0ENO(_d256), .FORW_UA0WEO(_d257), .FORW_LA0CLKO(_d258), .FORW_LA0ENO(_d259), .FORW_LA0WEO(_d260),
                   .FORW_UA1CLKO(_d261), .FORW_UA1ENO(_d262), .FORW_UA1WEO(_d263), .FORW_LA1CLKO(_d264), .FORW_LA1ENO(_d265), .FORW_LA1WEO(_d266),
                   .FORW_UB0CLKO(_d267), .FORW_UB0ENO(_d268), .FORW_UB0WEO(_d269), .FORW_LB0CLKO(_d270), .FORW_LB0ENO(_d271), .FORW_LB0WEO(_d272),
                   .FORW_UB1CLKO(_d273), .FORW_UB1ENO(_d274), .FORW_UB1WEO(_d275), .FORW_LB1CLKO(_d276), .FORW_LB1ENO(_d277), .FORW_LB1WEO(_d278),
                   .CLOCKA({_d279, _d280, _d281, _d282}),
                   .CLOCKB({_d283, _d284, _d285, _d286}),
                   .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .CLKB({1'b1, 1'b1, 1'b1, na411_9}),
                   .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .GLWEA({1'b1, 1'b1, 1'b1, na412_10}),
                   .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0({na415_10, na419_9, na421_10, na445_9, na447_10, na458_9, na459_10, na460_9, na461_10, na463_9, na468_10,
                  na471_9, na472_10, na473_9, na474_10, na481_9}),
                   .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB0({na482_10, na484_9, na485_10, na489_9, na490_10, na491_9, na492_10, na493_9, na494_10, na495_9, na496_10,
                  na497_9, na498_10, na499_9, na500_10, na501_9}),
                   .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .DIA({na502_10, na503_9, na504_10, na505_9, na506_10, na507_9, na508_10, na509_9, na510_10, na511_9, na512_10, na513_9,
                  na514_10, na515_9, na516_10, na517_9, na518_10, na519_9, na520_10, na521_9, na522_10, na523_9, na524_10, na525_9,
                  na526_10, na527_9, na528_10, na529_9, na530_10, na531_9, na532_10, na533_9, na534_10, na535_9, na536_10, na537_9,
                  na538_10, na539_9, na540_10, na541_9}),
                   .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEA({na542_10, na543_9, na544_10, na545_9, na546_10, na547_9, na548_10, na549_9, na550_10, na551_9, na552_10, na553_9,
                  na554_10, na555_9, na556_10, na557_9, na558_10, na559_9, na560_10, na561_9, na562_10, na563_9, na564_10, na565_9,
                  na566_10, na567_9, na568_10, na569_9, na570_10, na571_9, na572_10, na573_9, na574_10, na575_9, na576_10, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .CLOCK1(na250_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                   .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                   .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                   .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                   .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_01_04_05_00_60_00_0C_00_00_00_03_13_00_00_00_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a399 ( .DOA({_d287, _d288, _d289, _d290, _d291, _d292, _d293, _d294, _d295, _d296, _d297, _d298, _d299, _d300, _d301, _d302,
                  _d303, _d304, _d305, _d306, _d307, _d308, _d309, _d310, _d311, _d312, _d313, _d314, _d315, _d316, _d317, _d318, _d319,
                  _d320, _d321, _d322, _d323, _d324, _d325, _d326}),
                   .DOAX({_d327, _d328, _d329, _d330, _d331, _d332, _d333, _d334, _d335, _d336, _d337, _d338, _d339, _d340, _d341,
                  _d342, _d343, _d344, _d345, _d346, _d347, _d348, _d349, _d350, _d351, _d352, _d353, _d354, _d355, _d356, _d357, _d358,
                  _d359, _d360, _d361, _d362, _d363, _d364, _d365, _d366}),
                   .DOB({_d367, _d368, _d369, _d370, _d371, _d372, _d373, _d374, _d375, _d376, _d377, _d378, _d379, _d380, _d381, _d382,
                  _d383, _d384, _d385, _d386, _d387, _d388, _d389, _d390, _d391, _d392, _d393, _d394, _d395, _d396, _d397, _d398, _d399,
                  _d400, _d401, _d402, _d403, na399_118, na399_119, na399_120}),
                   .DOBX({_d404, _d405, _d406, _d407, _d408, _d409, _d410, _d411, _d412, _d413, _d414, _d415, _d416, _d417, _d418,
                  _d419, _d420, _d421, _d422, _d423, _d424, _d425, _d426, _d427, _d428, _d429, _d430, _d431, _d432, _d433, _d434, _d435,
                  _d436, _d437, _d438, _d439, _d440, _d441, _d442, _d443}),
                   .ECC1B_ERRA({_d444, _d445, _d446, _d447}),
                   .ECC1B_ERRB({_d448, _d449, _d450, _d451}),
                   .ECC2B_ERRA({_d452, _d453, _d454, _d455}),
                   .ECC2B_ERRB({_d456, _d457, _d458, _d459}),
                   .FORW_CAS_WRAO(_d460), .FORW_CAS_WRBO(_d461), .FORW_CAS_BMAO(_d462), .FORW_CAS_BMBO(_d463), .FORW_CAS_RDAO(_d464),
                   .FORW_CAS_RDBO(_d465), .FORW_UADDRAO({_d466, _d467, _d468, _d469, _d470, _d471, _d472, _d473, _d474, _d475, _d476,
                  _d477, _d478, _d479, _d480, _d481}),
                   .FORW_LADDRAO({_d482, _d483, _d484, _d485, _d486, _d487, _d488, _d489, _d490, _d491, _d492, _d493, _d494, _d495,
                  _d496, _d497}),
                   .FORW_UADDRBO({_d498, _d499, _d500, _d501, _d502, _d503, _d504, _d505, _d506, _d507, _d508, _d509, _d510, _d511,
                  _d512, _d513}),
                   .FORW_LADDRBO({_d514, _d515, _d516, _d517, _d518, _d519, _d520, _d521, _d522, _d523, _d524, _d525, _d526, _d527,
                  _d528, _d529}),
                   .FORW_UA0CLKO(_d530), .FORW_UA0ENO(_d531), .FORW_UA0WEO(_d532), .FORW_LA0CLKO(_d533), .FORW_LA0ENO(_d534), .FORW_LA0WEO(_d535),
                   .FORW_UA1CLKO(_d536), .FORW_UA1ENO(_d537), .FORW_UA1WEO(_d538), .FORW_LA1CLKO(_d539), .FORW_LA1ENO(_d540), .FORW_LA1WEO(_d541),
                   .FORW_UB0CLKO(_d542), .FORW_UB0ENO(_d543), .FORW_UB0WEO(_d544), .FORW_LB0CLKO(_d545), .FORW_LB0ENO(_d546), .FORW_LB0WEO(_d547),
                   .FORW_UB1CLKO(_d548), .FORW_UB1ENO(_d549), .FORW_UB1WEO(_d550), .FORW_LB1CLKO(_d551), .FORW_LB1ENO(_d552), .FORW_LB1WEO(_d553),
                   .CLOCKA({_d554, _d555, _d556, _d557}),
                   .CLOCKB({_d558, _d559, _d560, _d561}),
                   .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .CLKB({1'b1, 1'b1, 1'b1, na580_9}),
                   .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .GLWEA({1'b1, 1'b1, 1'b1, na581_10}),
                   .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0({na582_10, na583_9, na584_10, na585_9, na586_10, na587_9, na588_10, na589_9, na590_10, na591_9, na592_10,
                  na593_9, na594_10, na595_9, na596_10, na597_9}),
                   .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB0({na598_10, na599_9, na600_10, na601_9, na602_10, na603_9, na604_10, na605_9, na606_10, na607_9, na608_10,
                  na609_9, na610_10, na611_9, na612_10, na613_9}),
                   .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .DIA({na614_10, na615_9, na616_10, na617_9, na618_10, na619_9, na620_10, na621_9, na622_10, na623_9, na624_10, na625_9,
                  na626_10, na627_9, na628_10, na629_9, na630_10, na631_9, na632_10, na633_9, na634_10, na635_9, na636_10, na637_9,
                  na638_10, na639_9, na640_10, na641_9, na642_10, na643_9, na644_10, na645_9, na646_10, na647_9, na648_10, na649_9,
                  na650_10, na651_9, na652_10, na653_9}),
                   .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEA({na654_10, na655_9, na656_10, na657_9, na658_10, na659_9, na660_10, na661_9, na662_10, na663_9, na664_10, na665_9,
                  na666_10, na667_9, na668_10, na669_9, na670_10, na671_9, na672_10, na673_9, na674_10, na675_9, na676_10, na677_9,
                  na678_10, na679_9, na680_10, na681_9, na682_10, na683_9, na684_10, na685_9, na686_10, na687_9, na688_10, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .CLOCK1(na250_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                   .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                   .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                   .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                   .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_01_04_05_00_60_00_0C_00_00_00_03_13_00_00_00_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a400 ( .DOA({_d562, _d563, _d564, _d565, _d566, _d567, _d568, _d569, _d570, _d571, _d572, _d573, _d574, _d575, _d576, _d577,
                  _d578, _d579, _d580, _d581, _d582, _d583, _d584, _d585, _d586, _d587, _d588, _d589, _d590, _d591, _d592, _d593, _d594,
                  _d595, _d596, _d597, _d598, _d599, _d600, _d601}),
                   .DOAX({_d602, _d603, _d604, _d605, _d606, _d607, _d608, _d609, _d610, _d611, _d612, _d613, _d614, _d615, _d616,
                  _d617, _d618, _d619, _d620, _d621, _d622, _d623, _d624, _d625, _d626, _d627, _d628, _d629, _d630, _d631, _d632, _d633,
                  _d634, _d635, _d636, _d637, _d638, _d639, _d640, _d641}),
                   .DOB({_d642, _d643, _d644, _d645, _d646, _d647, _d648, _d649, _d650, _d651, _d652, _d653, _d654, _d655, _d656, _d657,
                  _d658, _d659, _d660, _d661, _d662, _d663, _d664, _d665, _d666, _d667, _d668, _d669, _d670, _d671, _d672, _d673, _d674,
                  _d675, _d676, _d677, _d678, na400_118, na400_119, na400_120}),
                   .DOBX({_d679, _d680, _d681, _d682, _d683, _d684, _d685, _d686, _d687, _d688, _d689, _d690, _d691, _d692, _d693,
                  _d694, _d695, _d696, _d697, _d698, _d699, _d700, _d701, _d702, _d703, _d704, _d705, _d706, _d707, _d708, _d709, _d710,
                  _d711, _d712, _d713, _d714, _d715, _d716, _d717, _d718}),
                   .ECC1B_ERRA({_d719, _d720, _d721, _d722}),
                   .ECC1B_ERRB({_d723, _d724, _d725, _d726}),
                   .ECC2B_ERRA({_d727, _d728, _d729, _d730}),
                   .ECC2B_ERRB({_d731, _d732, _d733, _d734}),
                   .FORW_CAS_WRAO(_d735), .FORW_CAS_WRBO(_d736), .FORW_CAS_BMAO(_d737), .FORW_CAS_BMBO(_d738), .FORW_CAS_RDAO(_d739),
                   .FORW_CAS_RDBO(_d740), .FORW_UADDRAO({_d741, _d742, _d743, _d744, _d745, _d746, _d747, _d748, _d749, _d750, _d751,
                  _d752, _d753, _d754, _d755, _d756}),
                   .FORW_LADDRAO({_d757, _d758, _d759, _d760, _d761, _d762, _d763, _d764, _d765, _d766, _d767, _d768, _d769, _d770,
                  _d771, _d772}),
                   .FORW_UADDRBO({_d773, _d774, _d775, _d776, _d777, _d778, _d779, _d780, _d781, _d782, _d783, _d784, _d785, _d786,
                  _d787, _d788}),
                   .FORW_LADDRBO({_d789, _d790, _d791, _d792, _d793, _d794, _d795, _d796, _d797, _d798, _d799, _d800, _d801, _d802,
                  _d803, _d804}),
                   .FORW_UA0CLKO(_d805), .FORW_UA0ENO(_d806), .FORW_UA0WEO(_d807), .FORW_LA0CLKO(_d808), .FORW_LA0ENO(_d809), .FORW_LA0WEO(_d810),
                   .FORW_UA1CLKO(_d811), .FORW_UA1ENO(_d812), .FORW_UA1WEO(_d813), .FORW_LA1CLKO(_d814), .FORW_LA1ENO(_d815), .FORW_LA1WEO(_d816),
                   .FORW_UB0CLKO(_d817), .FORW_UB0ENO(_d818), .FORW_UB0WEO(_d819), .FORW_LB0CLKO(_d820), .FORW_LB0ENO(_d821), .FORW_LB0WEO(_d822),
                   .FORW_UB1CLKO(_d823), .FORW_UB1ENO(_d824), .FORW_UB1WEO(_d825), .FORW_LB1CLKO(_d826), .FORW_LB1ENO(_d827), .FORW_LB1WEO(_d828),
                   .CLOCKA({_d829, _d830, _d831, _d832}),
                   .CLOCKB({_d833, _d834, _d835, _d836}),
                   .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .CLKB({1'b1, 1'b1, 1'b1, na692_9}),
                   .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .GLWEA({1'b1, 1'b1, 1'b1, na693_10}),
                   .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0({na694_10, na695_9, na696_10, na697_9, na698_10, na699_9, na700_10, na701_9, na702_10, na703_9, na704_10,
                  na705_9, na706_10, na707_9, na708_10, na709_9}),
                   .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB0({na710_10, na711_9, na712_10, na713_9, na714_10, na715_9, na716_10, na717_9, na718_10, na719_9, na720_10,
                  na721_9, na722_10, na723_9, na724_10, na725_9}),
                   .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .DIA({na726_10, na727_9, na728_10, na729_9, na730_10, na731_9, na732_10, na733_9, na734_10, na735_9, na736_10, na737_9,
                  na738_10, na739_9, na740_10, na741_9, na742_10, na743_9, na744_10, na745_9, na746_10, na747_9, na748_10, na749_9,
                  na750_10, na751_9, na752_10, na753_9, na754_10, na755_9, na756_10, na757_9, na758_10, na759_9, na760_10, na761_9,
                  na762_10, na763_9, na764_10, na765_9}),
                   .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEA({na766_10, na767_9, na768_10, na769_9, na770_10, na771_9, na772_10, na773_9, na774_10, na775_9, na776_10, na777_9,
                  na778_10, na779_9, na780_10, na781_9, na782_10, na783_9, na784_10, na785_9, na786_10, na787_9, na788_10, na789_9,
                  na790_10, na791_9, na792_10, na793_9, na794_10, na795_9, na796_10, na797_9, na798_10, na799_9, na800_10, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .CLOCK1(na250_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                   .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                   .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                   .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                   .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_01_04_05_00_60_00_0C_00_00_00_03_13_00_00_00_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a401 ( .DOA({_d837, _d838, _d839, _d840, _d841, _d842, _d843, _d844, _d845, _d846, _d847, _d848, _d849, _d850, _d851, _d852,
                  _d853, _d854, _d855, _d856, _d857, _d858, _d859, _d860, _d861, _d862, _d863, _d864, _d865, _d866, _d867, _d868, _d869,
                  _d870, _d871, _d872, _d873, _d874, _d875, _d876}),
                   .DOAX({_d877, _d878, _d879, _d880, _d881, _d882, _d883, _d884, _d885, _d886, _d887, _d888, _d889, _d890, _d891,
                  _d892, _d893, _d894, _d895, _d896, _d897, _d898, _d899, _d900, _d901, _d902, _d903, _d904, _d905, _d906, _d907, _d908,
                  _d909, _d910, _d911, _d912, _d913, _d914, _d915, _d916}),
                   .DOB({_d917, _d918, _d919, _d920, _d921, _d922, _d923, _d924, _d925, _d926, _d927, _d928, _d929, _d930, _d931, _d932,
                  _d933, _d934, _d935, _d936, _d937, _d938, _d939, _d940, _d941, _d942, _d943, _d944, _d945, _d946, _d947, _d948, _d949,
                  _d950, _d951, _d952, _d953, na401_118, na401_119, na401_120}),
                   .DOBX({_d954, _d955, _d956, _d957, _d958, _d959, _d960, _d961, _d962, _d963, _d964, _d965, _d966, _d967, _d968,
                  _d969, _d970, _d971, _d972, _d973, _d974, _d975, _d976, _d977, _d978, _d979, _d980, _d981, _d982, _d983, _d984, _d985,
                  _d986, _d987, _d988, _d989, _d990, _d991, _d992, _d993}),
                   .ECC1B_ERRA({_d994, _d995, _d996, _d997}),
                   .ECC1B_ERRB({_d998, _d999, _d1000, _d1001}),
                   .ECC2B_ERRA({_d1002, _d1003, _d1004, _d1005}),
                   .ECC2B_ERRB({_d1006, _d1007, _d1008, _d1009}),
                   .FORW_CAS_WRAO(_d1010), .FORW_CAS_WRBO(_d1011), .FORW_CAS_BMAO(_d1012), .FORW_CAS_BMBO(_d1013), .FORW_CAS_RDAO(_d1014),
                   .FORW_CAS_RDBO(_d1015), .FORW_UADDRAO({_d1016, _d1017, _d1018, _d1019, _d1020, _d1021, _d1022, _d1023, _d1024, _d1025,
                  _d1026, _d1027, _d1028, _d1029, _d1030, _d1031}),
                   .FORW_LADDRAO({_d1032, _d1033, _d1034, _d1035, _d1036, _d1037, _d1038, _d1039, _d1040, _d1041, _d1042, _d1043, _d1044,
                  _d1045, _d1046, _d1047}),
                   .FORW_UADDRBO({_d1048, _d1049, _d1050, _d1051, _d1052, _d1053, _d1054, _d1055, _d1056, _d1057, _d1058, _d1059, _d1060,
                  _d1061, _d1062, _d1063}),
                   .FORW_LADDRBO({_d1064, _d1065, _d1066, _d1067, _d1068, _d1069, _d1070, _d1071, _d1072, _d1073, _d1074, _d1075, _d1076,
                  _d1077, _d1078, _d1079}),
                   .FORW_UA0CLKO(_d1080), .FORW_UA0ENO(_d1081), .FORW_UA0WEO(_d1082), .FORW_LA0CLKO(_d1083), .FORW_LA0ENO(_d1084),
                   .FORW_LA0WEO(_d1085), .FORW_UA1CLKO(_d1086), .FORW_UA1ENO(_d1087), .FORW_UA1WEO(_d1088), .FORW_LA1CLKO(_d1089),
                   .FORW_LA1ENO(_d1090), .FORW_LA1WEO(_d1091), .FORW_UB0CLKO(_d1092), .FORW_UB0ENO(_d1093), .FORW_UB0WEO(_d1094), .FORW_LB0CLKO(_d1095),
                   .FORW_LB0ENO(_d1096), .FORW_LB0WEO(_d1097), .FORW_UB1CLKO(_d1098), .FORW_UB1ENO(_d1099), .FORW_UB1WEO(_d1100), .FORW_LB1CLKO(_d1101),
                   .FORW_LB1ENO(_d1102), .FORW_LB1WEO(_d1103), .CLOCKA({_d1104, _d1105, _d1106, _d1107}),
                   .CLOCKB({_d1108, _d1109, _d1110, _d1111}),
                   .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .CLKB({1'b1, 1'b1, 1'b1, na804_9}),
                   .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .GLWEA({1'b1, 1'b1, 1'b1, na805_10}),
                   .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0({na806_10, na807_9, na808_10, na809_9, na810_10, na811_9, na812_10, na813_9, na814_10, na815_9, na816_10,
                  na817_9, na818_10, na819_9, na820_10, na821_9}),
                   .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB0({na822_10, na823_9, na824_10, na825_9, na826_10, na827_9, na828_10, na829_9, na830_10, na831_9, na832_10,
                  na833_9, na834_10, na835_9, na836_10, na837_9}),
                   .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .DIA({na838_10, na839_9, na840_10, na841_9, na842_10, na843_9, na844_10, na845_9, na846_10, na847_9, na848_10, na849_9,
                  na850_10, na851_9, na852_10, na853_9, na854_10, na855_9, na856_10, na857_9, na858_10, na859_9, na860_10, na861_9,
                  na862_10, na863_9, na864_10, na865_9, na866_10, na867_9, na868_10, na869_9, na870_10, na871_9, na872_10, na873_9,
                  na874_10, na875_9, na876_10, na877_9}),
                   .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEA({na878_10, na879_9, na880_10, na881_9, na882_10, na883_9, na884_10, na885_9, na886_10, na887_9, na888_10, na889_9,
                  na890_10, na891_9, na892_10, na893_9, na894_10, na895_9, na896_10, na897_9, na898_10, na899_9, na900_10, na901_9,
                  na902_10, na903_9, na904_10, na905_9, na906_10, na907_9, na908_10, na909_9, na910_10, na911_9, na912_10, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .CLOCK1(na250_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                   .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                   .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                   .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                   .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
CC_USR_RSTN            _a402 ( .USR_RSTN(na402_1) );
// C_/RAM_I1///      x45y128     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a403_2 ( .OUT(na403_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na396_4), .CP_O(1'b0) );
// C_MX2b////      x48y44     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a404_1 ( .OUT(na404_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na916_2), .IN5(1'b0), .IN6(na920_2), .IN7(1'b0), .IN8(na220_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x36y39     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a405_1 ( .OUT(na405_1), .IN1(1'b1), .IN2(na1_1), .IN3(1'b0), .IN4(1'b0), .IN5(na73_2), .IN6(na8_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x41y39     80'h00_0060_00_0000_0C0E_FF7A
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a406_4 ( .OUT(na406_2), .IN1(na11_2), .IN2(1'b0), .IN3(~na4_1), .IN4(~na12_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x51y35     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a407_2 ( .OUT(na407_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a407_6 ( .COUTY1(na407_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na407_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a408 ( .PCLK0(na408_1), .PCLK1(na408_2), .PCLK2(_d1112), .PCLK3(_d1113), .CLK0(na390_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0),
                   .SER_CLK(1'b0), .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_////RAM_I2      x1y66     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a409_5 ( .OUT(na409_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na402_1), .CP_O(1'b0) );
// C_///AND/      x36y43     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a410_4 ( .OUT(na410_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na156_2), .IN4(na30_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y49     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a411_1 ( .OUT(na411_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na392_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a411_6 ( .RAM_O1(na411_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na411_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x27y49     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a412_4 ( .OUT(na412_2), .IN1(1'b1), .IN2(na150_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a412_6 ( .RAM_O2(na412_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na412_2), .COMP_OUT(1'b0) );
// C_MX2b////      x37y43     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a413_1 ( .OUT(na413_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na916_2), .IN5(na73_1), .IN6(1'b0), .IN7(na15_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x42y40     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a414_1 ( .OUT(na414_1), .IN1(1'b1), .IN2(~na1_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na15_2), .IN8(na87_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y56     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a415_4 ( .OUT(na415_2), .IN1(1'b1), .IN2(na97_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a415_6 ( .RAM_O2(na415_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na415_2), .COMP_OUT(1'b0) );
// C_MX2b////      x35y51     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a416_1 ( .OUT(na416_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na22_1), .IN5(1'b0), .IN6(na121_1), .IN7(1'b0), .IN8(na21_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x30y43     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a417_1 ( .OUT(na417_1), .IN1(na24_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na23_1), .IN6(na121_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x34y37     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a418_1 ( .OUT(na418_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na84_2), .IN6(1'b0), .IN7(na40_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y56     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a419_1 ( .OUT(na419_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na97_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a419_6 ( .RAM_O1(na419_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na419_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x45y37     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a420_1 ( .OUT(na420_1), .IN1(1'b1), .IN2(~na1_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na118_2), .IN8(na226_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y55     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a421_4 ( .OUT(na421_2), .IN1(1'b1), .IN2(na99_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a421_6 ( .RAM_O2(na421_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na421_2), .COMP_OUT(1'b0) );
// C_MX2b////      x49y42     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a422_1 ( .OUT(na422_1), .IN1(1'b1), .IN2(na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na32_1), .IN6(na247_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x42y42     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a423_1 ( .OUT(na423_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na162_2), .IN7(na156_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y43     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a424_1 ( .OUT(na424_1), .IN1(1'b1), .IN2(na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na38_1), .IN6(na237_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y42     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a425_1 ( .OUT(na425_1), .IN1(1'b1), .IN2(~na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na235_2), .IN6(na39_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x44y40     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a426_1 ( .OUT(na426_1), .IN1(1'b1), .IN2(~na1_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na40_1), .IN8(na230_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y37     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a427_1 ( .OUT(na427_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na41_1), .IN6(1'b0), .IN7(na232_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x45y45     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a428_1 ( .OUT(na428_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na19_2), .IN6(1'b0), .IN7(na232_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x46y43     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a429_1 ( .OUT(na429_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na916_2), .IN5(1'b0), .IN6(na921_2), .IN7(1'b0), .IN8(na220_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x42y37     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a430_1 ( .OUT(na430_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na64_2), .IN6(1'b0), .IN7(na228_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x43y35     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a431_1 ( .OUT(na431_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na64_1), .IN6(1'b0), .IN7(na228_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x34y41     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a432_1 ( .OUT(na432_1), .IN1(1'b1), .IN2(na1_1), .IN3(1'b0), .IN4(1'b0), .IN5(na64_2), .IN6(na102_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y41     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a433_1 ( .OUT(na433_1), .IN1(1'b1), .IN2(na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na32_2), .IN6(na247_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y39     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a434_1 ( .OUT(na434_1), .IN1(1'b1), .IN2(~na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na235_1), .IN6(na69_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y37     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a435_1 ( .OUT(na435_1), .IN1(1'b1), .IN2(~na1_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na40_2), .IN8(na230_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x41y40     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a436_1 ( .OUT(na436_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na117_2), .IN6(1'b0), .IN7(na118_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y45     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a437_1 ( .OUT(na437_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na73_1), .IN6(1'b0), .IN7(na224_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x44y38     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a438_1 ( .OUT(na438_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na73_2), .IN6(1'b0), .IN7(na224_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x36y34     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a439_1 ( .OUT(na439_1), .IN1(1'b1), .IN2(~na138_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na914_2), .IN8(~na955_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x48y46     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a440_1 ( .OUT(na440_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na79_1), .IN6(1'b0), .IN7(na222_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y35     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a441_1 ( .OUT(na441_1), .IN1(1'b1), .IN2(~na138_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na959_2), .IN8(~na689_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x33y37     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a442_1 ( .OUT(na442_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na84_1), .IN6(1'b0), .IN7(na40_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y40     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a443_1 ( .OUT(na443_1), .IN1(1'b1), .IN2(na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na85_1), .IN6(na239_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y38     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a444_1 ( .OUT(na444_1), .IN1(1'b1), .IN2(na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na85_2), .IN6(na239_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y55     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a445_1 ( .OUT(na445_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na99_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a445_6 ( .RAM_O1(na445_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na445_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x43y37     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a446_1 ( .OUT(na446_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na916_2), .IN5(na79_1), .IN6(1'b0), .IN7(na91_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y54     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a447_4 ( .OUT(na447_2), .IN1(na84_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a447_6 ( .RAM_O2(na447_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na447_2), .COMP_OUT(1'b0) );
// C_MX2b////      x49y35     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a448_1 ( .OUT(na448_1), .IN1(1'b1), .IN2(~na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na241_2), .IN6(na94_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y42     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a449_1 ( .OUT(na449_1), .IN1(1'b1), .IN2(na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na100_2), .IN6(na243_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x41y38     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a450_1 ( .OUT(na450_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na916_2), .IN5(na79_2), .IN6(1'b0), .IN7(na91_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x33y41     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a451_1 ( .OUT(na451_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na916_2), .IN5(1'b0), .IN6(na97_1), .IN7(1'b0), .IN8(na6_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y45     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a452_1 ( .OUT(na452_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na916_2), .IN5(1'b0), .IN6(na97_2), .IN7(1'b0), .IN8(na6_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x33y40     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a453_1 ( .OUT(na453_1), .IN1(1'b1), .IN2(na1_1), .IN3(1'b0), .IN4(1'b0), .IN5(na19_2), .IN6(na99_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y37     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a454_1 ( .OUT(na454_1), .IN1(1'b1), .IN2(na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na100_1), .IN6(na243_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y38     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a455_1 ( .OUT(na455_1), .IN1(1'b1), .IN2(~na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na245_1), .IN6(na141_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x34y38     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a456_1 ( .OUT(na456_1), .IN1(1'b1), .IN2(na1_1), .IN3(1'b0), .IN4(1'b0), .IN5(na64_1), .IN6(na102_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x39y37     80'h00_0018_00_0000_0888_CBCD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a457_1 ( .OUT(na457_1), .IN1(~na25_1), .IN2(na1_1), .IN3(1'b0), .IN4(na7_2), .IN5(na939_2), .IN6(~na1_1), .IN7(1'b0), .IN8(na7_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y54     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a458_1 ( .OUT(na458_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na84_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a458_6 ( .RAM_O1(na458_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na458_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y53     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a459_4 ( .OUT(na459_2), .IN1(1'b1), .IN2(na102_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a459_6 ( .RAM_O2(na459_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na459_2), .COMP_OUT(1'b0) );
// C_AND////      x28y53     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a460_1 ( .OUT(na460_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na102_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a460_6 ( .RAM_O1(na460_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na460_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y52     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a461_4 ( .OUT(na461_2), .IN1(na117_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a461_6 ( .RAM_O2(na461_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na461_2), .COMP_OUT(1'b0) );
// C_MX2b////      x40y50     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a462_1 ( .OUT(na462_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na22_1), .IN5(na5_1), .IN6(1'b0), .IN7(na107_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y52     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a463_1 ( .OUT(na463_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na117_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a463_6 ( .RAM_O1(na463_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na463_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x38y50     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a464_1 ( .OUT(na464_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3_1), .IN6(1'b1), .IN7(1'b1), .IN8(na30_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x29y44     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a465_1 ( .OUT(na465_1), .IN1(~na24_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na5_1), .IN6(na935_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x39y51     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a466_1 ( .OUT(na466_1), .IN1(~na24_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na120_1), .IN8(na936_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x38y52     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a467_1 ( .OUT(na467_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3_1), .IN6(na114_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y51     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a468_4 ( .OUT(na468_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a468_6 ( .RAM_O2(na468_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na468_2), .COMP_OUT(1'b0) );
// C_MX2b////      x41y37     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a469_1 ( .OUT(na469_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na117_1), .IN6(1'b0), .IN7(na118_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x45y44     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a470_1 ( .OUT(na470_1), .IN1(1'b1), .IN2(~na1_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na118_1), .IN8(na226_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y51     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a471_1 ( .OUT(na471_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na8_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a471_6 ( .RAM_O1(na471_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na471_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y50     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a472_4 ( .OUT(na472_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a472_6 ( .RAM_O2(na472_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na472_2), .COMP_OUT(1'b0) );
// C_AND////      x28y50     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a473_1 ( .OUT(na473_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a473_6 ( .RAM_O1(na473_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na473_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y49     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a474_4 ( .OUT(na474_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a474_6 ( .RAM_O2(na474_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na474_2), .COMP_OUT(1'b0) );
// C_MX2b////      x36y37     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a475_1 ( .OUT(na475_1), .IN1(1'b1), .IN2(na1_1), .IN3(1'b0), .IN4(1'b0), .IN5(na41_1), .IN6(na99_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y40     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a476_1 ( .OUT(na476_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na17_1), .IN5(1'b0), .IN6(na237_2), .IN7(1'b0), .IN8(na938_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y37     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a477_1 ( .OUT(na477_1), .IN1(1'b1), .IN2(~na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na245_2), .IN6(na141_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x45y38     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a478_1 ( .OUT(na478_1), .IN1(1'b1), .IN2(~na926_2), .IN3(1'b0), .IN4(1'b0), .IN5(na241_1), .IN6(na94_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x47y43     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a479_1 ( .OUT(na479_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na916_2), .IN5(na79_2), .IN6(1'b0), .IN7(na222_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y34     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a480_1 ( .OUT(na480_1), .IN1(1'b1), .IN2(~na138_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na915_1), .IN8(~na956_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a481_1 ( .OUT(na481_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a481_6 ( .RAM_O1(na481_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na481_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y56     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a482_4 ( .OUT(na482_2), .IN1(1'b1), .IN2(na136_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a482_6 ( .RAM_O2(na482_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na482_2), .COMP_OUT(1'b0) );
// C_///AND/      x41y46     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a483_4 ( .OUT(na483_2), .IN1(na153_1), .IN2(1'b1), .IN3(na27_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y56     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a484_1 ( .OUT(na484_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na135_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a484_6 ( .RAM_O1(na484_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na484_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y55     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a485_4 ( .OUT(na485_2), .IN1(na134_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a485_6 ( .RAM_O2(na485_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na485_2), .COMP_OUT(1'b0) );
// C_AND////      x41y47     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a486_1 ( .OUT(na486_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na939_2), .IN6(1'b1), .IN7(~na156_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x107y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a487_4 ( .OUT(na487_2), .IN1(1'b1), .IN2(1'b1), .IN3(na47_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a487_6 ( .RAM_O2(na487_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na487_2), .COMP_OUT(1'b0) );
// C_///AND/      x19y1     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a488_4 ( .OUT(na488_2), .IN1(1'b1), .IN2(1'b1), .IN3(na103_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a488_6 ( .RAM_O2(na488_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na488_2), .COMP_OUT(1'b0) );
// C_AND////      x37y55     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a489_1 ( .OUT(na489_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na133_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a489_6 ( .RAM_O1(na489_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na489_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y54     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a490_4 ( .OUT(na490_2), .IN1(1'b1), .IN2(na132_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a490_6 ( .RAM_O2(na490_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na490_2), .COMP_OUT(1'b0) );
// C_AND////      x37y54     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a491_1 ( .OUT(na491_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na131_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a491_6 ( .RAM_O1(na491_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na491_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y53     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a492_4 ( .OUT(na492_2), .IN1(1'b1), .IN2(1'b1), .IN3(na130_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a492_6 ( .RAM_O2(na492_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na492_2), .COMP_OUT(1'b0) );
// C_AND////      x37y53     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a493_1 ( .OUT(na493_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na129_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a493_6 ( .RAM_O1(na493_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na493_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y52     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a494_4 ( .OUT(na494_2), .IN1(1'b1), .IN2(na128_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a494_6 ( .RAM_O2(na494_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na494_2), .COMP_OUT(1'b0) );
// C_AND////      x37y52     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a495_1 ( .OUT(na495_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na127_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a495_6 ( .RAM_O1(na495_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na495_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y51     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a496_4 ( .OUT(na496_2), .IN1(1'b1), .IN2(na126_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a496_6 ( .RAM_O2(na496_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na496_2), .COMP_OUT(1'b0) );
// C_AND////      x37y51     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a497_1 ( .OUT(na497_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na125_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a497_6 ( .RAM_O1(na497_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na497_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y50     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a498_4 ( .OUT(na498_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na124_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a498_6 ( .RAM_O2(na498_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na498_2), .COMP_OUT(1'b0) );
// C_AND////      x37y50     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a499_1 ( .OUT(na499_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a499_6 ( .RAM_O1(na499_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na499_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y49     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a500_4 ( .OUT(na500_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a500_6 ( .RAM_O2(na500_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na500_2), .COMP_OUT(1'b0) );
// C_AND////      x37y49     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a501_1 ( .OUT(na501_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a501_6 ( .RAM_O1(na501_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na501_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a502_4 ( .OUT(na502_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a502_6 ( .RAM_O2(na502_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na502_2), .COMP_OUT(1'b0) );
// C_AND////      x30y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a503_1 ( .OUT(na503_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a503_6 ( .RAM_O1(na503_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na503_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a504_4 ( .OUT(na504_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a504_6 ( .RAM_O2(na504_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na504_2), .COMP_OUT(1'b0) );
// C_AND////      x30y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a505_1 ( .OUT(na505_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a505_6 ( .RAM_O1(na505_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na505_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a506_4 ( .OUT(na506_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a506_6 ( .RAM_O2(na506_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na506_2), .COMP_OUT(1'b0) );
// C_AND////      x32y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a507_1 ( .OUT(na507_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a507_6 ( .RAM_O1(na507_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na507_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a508_4 ( .OUT(na508_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a508_6 ( .RAM_O2(na508_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na508_2), .COMP_OUT(1'b0) );
// C_AND////      x32y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a509_1 ( .OUT(na509_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a509_6 ( .RAM_O1(na509_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na509_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y62     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a510_4 ( .OUT(na510_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a510_6 ( .RAM_O2(na510_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na510_2), .COMP_OUT(1'b0) );
// C_AND////      x32y62     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a511_1 ( .OUT(na511_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a511_6 ( .RAM_O1(na511_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na511_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y61     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a512_4 ( .OUT(na512_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a512_6 ( .RAM_O2(na512_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na512_2), .COMP_OUT(1'b0) );
// C_AND////      x32y61     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a513_1 ( .OUT(na513_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a513_6 ( .RAM_O1(na513_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na513_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y60     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a514_4 ( .OUT(na514_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a514_6 ( .RAM_O2(na514_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na514_2), .COMP_OUT(1'b0) );
// C_AND////      x32y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a515_1 ( .OUT(na515_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a515_6 ( .RAM_O1(na515_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na515_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y59     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a516_4 ( .OUT(na516_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a516_6 ( .RAM_O2(na516_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na516_2), .COMP_OUT(1'b0) );
// C_AND////      x32y59     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a517_1 ( .OUT(na517_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a517_6 ( .RAM_O1(na517_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na517_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y58     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a518_4 ( .OUT(na518_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a518_6 ( .RAM_O2(na518_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na518_2), .COMP_OUT(1'b0) );
// C_AND////      x32y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a519_1 ( .OUT(na519_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a519_6 ( .RAM_O1(na519_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na519_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a520_4 ( .OUT(na520_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a520_6 ( .RAM_O2(na520_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na520_2), .COMP_OUT(1'b0) );
// C_AND////      x32y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a521_1 ( .OUT(na521_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a521_6 ( .RAM_O1(na521_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na521_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y56     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a522_4 ( .OUT(na522_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a522_6 ( .RAM_O2(na522_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na522_2), .COMP_OUT(1'b0) );
// C_AND////      x30y56     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a523_1 ( .OUT(na523_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a523_6 ( .RAM_O1(na523_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na523_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y55     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a524_4 ( .OUT(na524_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a524_6 ( .RAM_O2(na524_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na524_2), .COMP_OUT(1'b0) );
// C_AND////      x30y55     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a525_1 ( .OUT(na525_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a525_6 ( .RAM_O1(na525_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na525_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y56     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a526_4 ( .OUT(na526_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a526_6 ( .RAM_O2(na526_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na526_2), .COMP_OUT(1'b0) );
// C_AND////      x32y56     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a527_1 ( .OUT(na527_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a527_6 ( .RAM_O1(na527_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na527_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y55     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a528_4 ( .OUT(na528_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a528_6 ( .RAM_O2(na528_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na528_2), .COMP_OUT(1'b0) );
// C_AND////      x32y55     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a529_1 ( .OUT(na529_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a529_6 ( .RAM_O1(na529_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na529_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y54     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a530_4 ( .OUT(na530_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a530_6 ( .RAM_O2(na530_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na530_2), .COMP_OUT(1'b0) );
// C_AND////      x32y54     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a531_1 ( .OUT(na531_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a531_6 ( .RAM_O1(na531_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na531_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y53     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a532_4 ( .OUT(na532_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a532_6 ( .RAM_O2(na532_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na532_2), .COMP_OUT(1'b0) );
// C_AND////      x32y53     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a533_1 ( .OUT(na533_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a533_6 ( .RAM_O1(na533_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na533_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y52     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a534_4 ( .OUT(na534_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a534_6 ( .RAM_O2(na534_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na534_2), .COMP_OUT(1'b0) );
// C_AND////      x32y52     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a535_1 ( .OUT(na535_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a535_6 ( .RAM_O1(na535_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na535_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y51     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a536_4 ( .OUT(na536_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a536_6 ( .RAM_O2(na536_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na536_2), .COMP_OUT(1'b0) );
// C_AND////      x32y51     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a537_1 ( .OUT(na537_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a537_6 ( .RAM_O1(na537_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na537_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y50     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a538_4 ( .OUT(na538_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a538_6 ( .RAM_O2(na538_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na538_2), .COMP_OUT(1'b0) );
// C_AND////      x32y50     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a539_1 ( .OUT(na539_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na390_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a539_6 ( .RAM_O1(na539_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na539_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y49     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a540_4 ( .OUT(na540_2), .IN1(1'b1), .IN2(na250_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a540_6 ( .RAM_O2(na540_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na540_2), .COMP_OUT(1'b0) );
// C_AND////      x32y49     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a541_1 ( .OUT(na541_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na403_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a541_6 ( .RAM_O1(na541_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na541_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a542_4 ( .OUT(na542_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a542_6 ( .RAM_O2(na542_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na542_2), .COMP_OUT(1'b0) );
// C_AND////      x29y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a543_1 ( .OUT(na543_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a543_6 ( .RAM_O1(na543_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na543_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a544_4 ( .OUT(na544_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a544_6 ( .RAM_O2(na544_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na544_2), .COMP_OUT(1'b0) );
// C_AND////      x29y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a545_1 ( .OUT(na545_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a545_6 ( .RAM_O1(na545_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na545_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a546_4 ( .OUT(na546_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a546_6 ( .RAM_O2(na546_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na546_2), .COMP_OUT(1'b0) );
// C_AND////      x31y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a547_1 ( .OUT(na547_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a547_6 ( .RAM_O1(na547_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na547_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a548_4 ( .OUT(na548_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a548_6 ( .RAM_O2(na548_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na548_2), .COMP_OUT(1'b0) );
// C_AND////      x31y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a549_1 ( .OUT(na549_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a549_6 ( .RAM_O1(na549_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na549_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y62     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a550_4 ( .OUT(na550_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a550_6 ( .RAM_O2(na550_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na550_2), .COMP_OUT(1'b0) );
// C_AND////      x31y62     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a551_1 ( .OUT(na551_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a551_6 ( .RAM_O1(na551_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na551_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y61     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a552_4 ( .OUT(na552_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a552_6 ( .RAM_O2(na552_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na552_2), .COMP_OUT(1'b0) );
// C_AND////      x31y61     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a553_1 ( .OUT(na553_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a553_6 ( .RAM_O1(na553_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na553_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y60     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a554_4 ( .OUT(na554_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a554_6 ( .RAM_O2(na554_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na554_2), .COMP_OUT(1'b0) );
// C_AND////      x31y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a555_1 ( .OUT(na555_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a555_6 ( .RAM_O1(na555_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na555_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y59     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a556_4 ( .OUT(na556_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a556_6 ( .RAM_O2(na556_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na556_2), .COMP_OUT(1'b0) );
// C_AND////      x31y59     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a557_1 ( .OUT(na557_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a557_6 ( .RAM_O1(na557_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na557_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y58     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a558_4 ( .OUT(na558_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a558_6 ( .RAM_O2(na558_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na558_2), .COMP_OUT(1'b0) );
// C_AND////      x31y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a559_1 ( .OUT(na559_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a559_6 ( .RAM_O1(na559_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na559_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a560_4 ( .OUT(na560_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a560_6 ( .RAM_O2(na560_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na560_2), .COMP_OUT(1'b0) );
// C_AND////      x31y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a561_1 ( .OUT(na561_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a561_6 ( .RAM_O1(na561_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na561_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y56     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a562_4 ( .OUT(na562_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a562_6 ( .RAM_O2(na562_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na562_2), .COMP_OUT(1'b0) );
// C_AND////      x29y56     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a563_1 ( .OUT(na563_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a563_6 ( .RAM_O1(na563_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na563_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y55     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a564_4 ( .OUT(na564_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a564_6 ( .RAM_O2(na564_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na564_2), .COMP_OUT(1'b0) );
// C_AND////      x29y55     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a565_1 ( .OUT(na565_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a565_6 ( .RAM_O1(na565_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na565_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y56     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a566_4 ( .OUT(na566_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a566_6 ( .RAM_O2(na566_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na566_2), .COMP_OUT(1'b0) );
// C_AND////      x31y56     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a567_1 ( .OUT(na567_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a567_6 ( .RAM_O1(na567_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na567_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y55     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a568_4 ( .OUT(na568_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a568_6 ( .RAM_O2(na568_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na568_2), .COMP_OUT(1'b0) );
// C_AND////      x31y55     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a569_1 ( .OUT(na569_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a569_6 ( .RAM_O1(na569_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na569_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y54     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a570_4 ( .OUT(na570_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a570_6 ( .RAM_O2(na570_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na570_2), .COMP_OUT(1'b0) );
// C_AND////      x31y54     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a571_1 ( .OUT(na571_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a571_6 ( .RAM_O1(na571_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na571_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y53     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a572_4 ( .OUT(na572_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a572_6 ( .RAM_O2(na572_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na572_2), .COMP_OUT(1'b0) );
// C_AND////      x31y53     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a573_1 ( .OUT(na573_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a573_6 ( .RAM_O1(na573_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na573_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y52     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a574_4 ( .OUT(na574_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a574_6 ( .RAM_O2(na574_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na574_2), .COMP_OUT(1'b0) );
// C_AND////      x31y52     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a575_1 ( .OUT(na575_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a575_6 ( .RAM_O1(na575_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na575_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y51     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a576_4 ( .OUT(na576_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a576_6 ( .RAM_O2(na576_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na576_2), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x34y50     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a577_2 ( .OUT(na577_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na398_118), .CP_O(1'b0) );
// C_////RAM_I2      x34y49     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a578_5 ( .OUT(na578_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na398_119), .CP_O(1'b0) );
// C_/RAM_I1///      x34y49     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a579_2 ( .OUT(na579_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na398_120), .CP_O(1'b0) );
// C_AND////      x35y33     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a580_1 ( .OUT(na580_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na392_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a580_6 ( .RAM_O1(na580_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na580_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x27y33     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a581_4 ( .OUT(na581_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na149_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a581_6 ( .RAM_O2(na581_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na581_2), .COMP_OUT(1'b0) );
// C_///AND/      x28y40     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a582_4 ( .OUT(na582_2), .IN1(1'b1), .IN2(na97_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a582_6 ( .RAM_O2(na582_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na582_2), .COMP_OUT(1'b0) );
// C_AND////      x28y40     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a583_1 ( .OUT(na583_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na97_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a583_6 ( .RAM_O1(na583_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na583_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y39     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a584_4 ( .OUT(na584_2), .IN1(1'b1), .IN2(na99_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a584_6 ( .RAM_O2(na584_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na584_2), .COMP_OUT(1'b0) );
// C_AND////      x28y39     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a585_1 ( .OUT(na585_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na99_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a585_6 ( .RAM_O1(na585_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na585_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y38     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a586_4 ( .OUT(na586_2), .IN1(na84_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a586_6 ( .RAM_O2(na586_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na586_2), .COMP_OUT(1'b0) );
// C_AND////      x28y38     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a587_1 ( .OUT(na587_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na84_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a587_6 ( .RAM_O1(na587_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na587_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y37     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a588_4 ( .OUT(na588_2), .IN1(1'b1), .IN2(na102_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a588_6 ( .RAM_O2(na588_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na588_2), .COMP_OUT(1'b0) );
// C_AND////      x28y37     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a589_1 ( .OUT(na589_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na102_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a589_6 ( .RAM_O1(na589_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na589_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y36     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a590_4 ( .OUT(na590_2), .IN1(na117_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a590_6 ( .RAM_O2(na590_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na590_2), .COMP_OUT(1'b0) );
// C_AND////      x28y36     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a591_1 ( .OUT(na591_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na117_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a591_6 ( .RAM_O1(na591_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na591_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y35     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a592_4 ( .OUT(na592_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a592_6 ( .RAM_O2(na592_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na592_2), .COMP_OUT(1'b0) );
// C_AND////      x28y35     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a593_1 ( .OUT(na593_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na8_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a593_6 ( .RAM_O1(na593_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na593_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y34     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a594_4 ( .OUT(na594_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a594_6 ( .RAM_O2(na594_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na594_2), .COMP_OUT(1'b0) );
// C_AND////      x28y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a595_1 ( .OUT(na595_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a595_6 ( .RAM_O1(na595_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na595_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a596_4 ( .OUT(na596_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a596_6 ( .RAM_O2(na596_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na596_2), .COMP_OUT(1'b0) );
// C_AND////      x28y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a597_1 ( .OUT(na597_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a597_6 ( .RAM_O1(na597_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na597_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y40     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a598_4 ( .OUT(na598_2), .IN1(1'b1), .IN2(na136_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a598_6 ( .RAM_O2(na598_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na598_2), .COMP_OUT(1'b0) );
// C_AND////      x37y40     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a599_1 ( .OUT(na599_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na135_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a599_6 ( .RAM_O1(na599_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na599_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y39     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a600_4 ( .OUT(na600_2), .IN1(na134_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a600_6 ( .RAM_O2(na600_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na600_2), .COMP_OUT(1'b0) );
// C_AND////      x37y39     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a601_1 ( .OUT(na601_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na133_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a601_6 ( .RAM_O1(na601_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na601_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y38     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a602_4 ( .OUT(na602_2), .IN1(1'b1), .IN2(na132_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a602_6 ( .RAM_O2(na602_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na602_2), .COMP_OUT(1'b0) );
// C_AND////      x37y38     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a603_1 ( .OUT(na603_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na131_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a603_6 ( .RAM_O1(na603_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na603_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y37     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a604_4 ( .OUT(na604_2), .IN1(1'b1), .IN2(1'b1), .IN3(na130_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a604_6 ( .RAM_O2(na604_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na604_2), .COMP_OUT(1'b0) );
// C_AND////      x37y37     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a605_1 ( .OUT(na605_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na129_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a605_6 ( .RAM_O1(na605_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na605_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y36     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a606_4 ( .OUT(na606_2), .IN1(1'b1), .IN2(na128_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a606_6 ( .RAM_O2(na606_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na606_2), .COMP_OUT(1'b0) );
// C_AND////      x37y36     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a607_1 ( .OUT(na607_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na127_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a607_6 ( .RAM_O1(na607_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na607_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y35     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a608_4 ( .OUT(na608_2), .IN1(1'b1), .IN2(na126_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a608_6 ( .RAM_O2(na608_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na608_2), .COMP_OUT(1'b0) );
// C_AND////      x37y35     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a609_1 ( .OUT(na609_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na125_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a609_6 ( .RAM_O1(na609_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na609_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y34     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a610_4 ( .OUT(na610_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na124_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a610_6 ( .RAM_O2(na610_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na610_2), .COMP_OUT(1'b0) );
// C_AND////      x37y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a611_1 ( .OUT(na611_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a611_6 ( .RAM_O1(na611_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na611_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a612_4 ( .OUT(na612_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a612_6 ( .RAM_O2(na612_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na612_2), .COMP_OUT(1'b0) );
// C_AND////      x37y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a613_1 ( .OUT(na613_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a613_6 ( .RAM_O1(na613_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na613_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a614_4 ( .OUT(na614_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a614_6 ( .RAM_O2(na614_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na614_2), .COMP_OUT(1'b0) );
// C_AND////      x30y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a615_1 ( .OUT(na615_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a615_6 ( .RAM_O1(na615_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na615_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a616_4 ( .OUT(na616_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a616_6 ( .RAM_O2(na616_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na616_2), .COMP_OUT(1'b0) );
// C_AND////      x30y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a617_1 ( .OUT(na617_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a617_6 ( .RAM_O1(na617_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na617_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a618_4 ( .OUT(na618_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a618_6 ( .RAM_O2(na618_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na618_2), .COMP_OUT(1'b0) );
// C_AND////      x32y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a619_1 ( .OUT(na619_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a619_6 ( .RAM_O1(na619_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na619_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a620_4 ( .OUT(na620_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a620_6 ( .RAM_O2(na620_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na620_2), .COMP_OUT(1'b0) );
// C_AND////      x32y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a621_1 ( .OUT(na621_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a621_6 ( .RAM_O1(na621_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na621_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y46     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a622_4 ( .OUT(na622_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a622_6 ( .RAM_O2(na622_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na622_2), .COMP_OUT(1'b0) );
// C_AND////      x32y46     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a623_1 ( .OUT(na623_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a623_6 ( .RAM_O1(na623_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na623_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y45     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a624_4 ( .OUT(na624_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a624_6 ( .RAM_O2(na624_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na624_2), .COMP_OUT(1'b0) );
// C_AND////      x32y45     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a625_1 ( .OUT(na625_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a625_6 ( .RAM_O1(na625_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na625_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y44     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a626_4 ( .OUT(na626_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a626_6 ( .RAM_O2(na626_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na626_2), .COMP_OUT(1'b0) );
// C_AND////      x32y44     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a627_1 ( .OUT(na627_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a627_6 ( .RAM_O1(na627_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na627_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y43     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a628_4 ( .OUT(na628_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a628_6 ( .RAM_O2(na628_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na628_2), .COMP_OUT(1'b0) );
// C_AND////      x32y43     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a629_1 ( .OUT(na629_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a629_6 ( .RAM_O1(na629_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na629_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y42     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a630_4 ( .OUT(na630_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a630_6 ( .RAM_O2(na630_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na630_2), .COMP_OUT(1'b0) );
// C_AND////      x32y42     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a631_1 ( .OUT(na631_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a631_6 ( .RAM_O1(na631_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na631_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y41     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a632_4 ( .OUT(na632_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a632_6 ( .RAM_O2(na632_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na632_2), .COMP_OUT(1'b0) );
// C_AND////      x32y41     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a633_1 ( .OUT(na633_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a633_6 ( .RAM_O1(na633_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na633_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a634_4 ( .OUT(na634_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a634_6 ( .RAM_O2(na634_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na634_2), .COMP_OUT(1'b0) );
// C_AND////      x30y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a635_1 ( .OUT(na635_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a635_6 ( .RAM_O1(na635_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na635_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a636_4 ( .OUT(na636_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a636_6 ( .RAM_O2(na636_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na636_2), .COMP_OUT(1'b0) );
// C_AND////      x30y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a637_1 ( .OUT(na637_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a637_6 ( .RAM_O1(na637_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na637_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a638_4 ( .OUT(na638_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a638_6 ( .RAM_O2(na638_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na638_2), .COMP_OUT(1'b0) );
// C_AND////      x32y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a639_1 ( .OUT(na639_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a639_6 ( .RAM_O1(na639_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na639_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a640_4 ( .OUT(na640_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a640_6 ( .RAM_O2(na640_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na640_2), .COMP_OUT(1'b0) );
// C_AND////      x32y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a641_1 ( .OUT(na641_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a641_6 ( .RAM_O1(na641_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na641_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y38     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a642_4 ( .OUT(na642_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a642_6 ( .RAM_O2(na642_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na642_2), .COMP_OUT(1'b0) );
// C_AND////      x32y38     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a643_1 ( .OUT(na643_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a643_6 ( .RAM_O1(na643_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na643_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y37     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a644_4 ( .OUT(na644_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a644_6 ( .RAM_O2(na644_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na644_2), .COMP_OUT(1'b0) );
// C_AND////      x32y37     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a645_1 ( .OUT(na645_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a645_6 ( .RAM_O1(na645_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na645_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y36     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a646_4 ( .OUT(na646_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a646_6 ( .RAM_O2(na646_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na646_2), .COMP_OUT(1'b0) );
// C_AND////      x32y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a647_1 ( .OUT(na647_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a647_6 ( .RAM_O1(na647_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na647_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y35     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a648_4 ( .OUT(na648_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a648_6 ( .RAM_O2(na648_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na648_2), .COMP_OUT(1'b0) );
// C_AND////      x32y35     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a649_1 ( .OUT(na649_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a649_6 ( .RAM_O1(na649_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na649_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y34     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a650_4 ( .OUT(na650_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a650_6 ( .RAM_O2(na650_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na650_2), .COMP_OUT(1'b0) );
// C_AND////      x32y34     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a651_1 ( .OUT(na651_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na390_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a651_6 ( .RAM_O1(na651_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na651_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y33     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a652_4 ( .OUT(na652_2), .IN1(1'b1), .IN2(na250_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a652_6 ( .RAM_O2(na652_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na652_2), .COMP_OUT(1'b0) );
// C_AND////      x32y33     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a653_1 ( .OUT(na653_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na403_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a653_6 ( .RAM_O1(na653_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na653_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a654_4 ( .OUT(na654_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a654_6 ( .RAM_O2(na654_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na654_2), .COMP_OUT(1'b0) );
// C_AND////      x29y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a655_1 ( .OUT(na655_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a655_6 ( .RAM_O1(na655_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na655_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a656_4 ( .OUT(na656_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a656_6 ( .RAM_O2(na656_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na656_2), .COMP_OUT(1'b0) );
// C_AND////      x29y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a657_1 ( .OUT(na657_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a657_6 ( .RAM_O1(na657_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na657_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a658_4 ( .OUT(na658_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a658_6 ( .RAM_O2(na658_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na658_2), .COMP_OUT(1'b0) );
// C_AND////      x31y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a659_1 ( .OUT(na659_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a659_6 ( .RAM_O1(na659_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na659_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a660_4 ( .OUT(na660_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a660_6 ( .RAM_O2(na660_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na660_2), .COMP_OUT(1'b0) );
// C_AND////      x31y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a661_1 ( .OUT(na661_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a661_6 ( .RAM_O1(na661_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na661_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y46     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a662_4 ( .OUT(na662_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a662_6 ( .RAM_O2(na662_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na662_2), .COMP_OUT(1'b0) );
// C_AND////      x31y46     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a663_1 ( .OUT(na663_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a663_6 ( .RAM_O1(na663_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na663_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y45     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a664_4 ( .OUT(na664_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a664_6 ( .RAM_O2(na664_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na664_2), .COMP_OUT(1'b0) );
// C_AND////      x31y45     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a665_1 ( .OUT(na665_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a665_6 ( .RAM_O1(na665_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na665_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y44     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a666_4 ( .OUT(na666_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a666_6 ( .RAM_O2(na666_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na666_2), .COMP_OUT(1'b0) );
// C_AND////      x31y44     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a667_1 ( .OUT(na667_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a667_6 ( .RAM_O1(na667_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na667_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y43     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a668_4 ( .OUT(na668_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a668_6 ( .RAM_O2(na668_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na668_2), .COMP_OUT(1'b0) );
// C_AND////      x31y43     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a669_1 ( .OUT(na669_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a669_6 ( .RAM_O1(na669_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na669_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y42     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a670_4 ( .OUT(na670_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a670_6 ( .RAM_O2(na670_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na670_2), .COMP_OUT(1'b0) );
// C_AND////      x31y42     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a671_1 ( .OUT(na671_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a671_6 ( .RAM_O1(na671_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na671_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y41     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a672_4 ( .OUT(na672_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a672_6 ( .RAM_O2(na672_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na672_2), .COMP_OUT(1'b0) );
// C_AND////      x31y41     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a673_1 ( .OUT(na673_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a673_6 ( .RAM_O1(na673_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na673_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a674_4 ( .OUT(na674_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a674_6 ( .RAM_O2(na674_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na674_2), .COMP_OUT(1'b0) );
// C_AND////      x29y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a675_1 ( .OUT(na675_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a675_6 ( .RAM_O1(na675_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na675_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a676_4 ( .OUT(na676_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a676_6 ( .RAM_O2(na676_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na676_2), .COMP_OUT(1'b0) );
// C_AND////      x29y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a677_1 ( .OUT(na677_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a677_6 ( .RAM_O1(na677_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na677_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a678_4 ( .OUT(na678_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a678_6 ( .RAM_O2(na678_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na678_2), .COMP_OUT(1'b0) );
// C_AND////      x31y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a679_1 ( .OUT(na679_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a679_6 ( .RAM_O1(na679_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na679_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a680_4 ( .OUT(na680_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a680_6 ( .RAM_O2(na680_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na680_2), .COMP_OUT(1'b0) );
// C_AND////      x31y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a681_1 ( .OUT(na681_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a681_6 ( .RAM_O1(na681_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na681_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y38     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a682_4 ( .OUT(na682_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a682_6 ( .RAM_O2(na682_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na682_2), .COMP_OUT(1'b0) );
// C_AND////      x31y38     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a683_1 ( .OUT(na683_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a683_6 ( .RAM_O1(na683_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na683_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y37     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a684_4 ( .OUT(na684_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a684_6 ( .RAM_O2(na684_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na684_2), .COMP_OUT(1'b0) );
// C_AND////      x31y37     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a685_1 ( .OUT(na685_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a685_6 ( .RAM_O1(na685_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na685_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y36     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a686_4 ( .OUT(na686_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a686_6 ( .RAM_O2(na686_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na686_2), .COMP_OUT(1'b0) );
// C_AND////      x31y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a687_1 ( .OUT(na687_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a687_6 ( .RAM_O1(na687_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na687_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y35     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a688_4 ( .OUT(na688_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a688_6 ( .RAM_O2(na688_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na688_2), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x34y34     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a689_2 ( .OUT(na689_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na399_118), .CP_O(1'b0) );
// C_////RAM_I2      x34y33     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a690_5 ( .OUT(na690_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na399_119), .CP_O(1'b0) );
// C_/RAM_I1///      x34y33     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a691_2 ( .OUT(na691_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na399_120), .CP_O(1'b0) );
// C_AND////      x35y65     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a692_1 ( .OUT(na692_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na392_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a692_6 ( .RAM_O1(na692_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na692_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x27y65     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a693_4 ( .OUT(na693_2), .IN1(1'b1), .IN2(1'b1), .IN3(na148_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a693_6 ( .RAM_O2(na693_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na693_2), .COMP_OUT(1'b0) );
// C_///AND/      x28y72     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a694_4 ( .OUT(na694_2), .IN1(1'b1), .IN2(na97_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a694_6 ( .RAM_O2(na694_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na694_2), .COMP_OUT(1'b0) );
// C_AND////      x28y72     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a695_1 ( .OUT(na695_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na97_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a695_6 ( .RAM_O1(na695_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na695_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y71     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a696_4 ( .OUT(na696_2), .IN1(1'b1), .IN2(na99_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a696_6 ( .RAM_O2(na696_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na696_2), .COMP_OUT(1'b0) );
// C_AND////      x28y71     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a697_1 ( .OUT(na697_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na99_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a697_6 ( .RAM_O1(na697_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na697_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y70     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a698_4 ( .OUT(na698_2), .IN1(na84_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a698_6 ( .RAM_O2(na698_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na698_2), .COMP_OUT(1'b0) );
// C_AND////      x28y70     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a699_1 ( .OUT(na699_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na84_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a699_6 ( .RAM_O1(na699_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na699_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y69     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a700_4 ( .OUT(na700_2), .IN1(1'b1), .IN2(na102_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a700_6 ( .RAM_O2(na700_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na700_2), .COMP_OUT(1'b0) );
// C_AND////      x28y69     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a701_1 ( .OUT(na701_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na102_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a701_6 ( .RAM_O1(na701_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na701_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y68     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a702_4 ( .OUT(na702_2), .IN1(na117_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a702_6 ( .RAM_O2(na702_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na702_2), .COMP_OUT(1'b0) );
// C_AND////      x28y68     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a703_1 ( .OUT(na703_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na117_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a703_6 ( .RAM_O1(na703_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na703_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y67     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a704_4 ( .OUT(na704_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a704_6 ( .RAM_O2(na704_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na704_2), .COMP_OUT(1'b0) );
// C_AND////      x28y67     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a705_1 ( .OUT(na705_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na8_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a705_6 ( .RAM_O1(na705_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na705_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y66     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a706_4 ( .OUT(na706_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a706_6 ( .RAM_O2(na706_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na706_2), .COMP_OUT(1'b0) );
// C_AND////      x28y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a707_1 ( .OUT(na707_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a707_6 ( .RAM_O1(na707_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na707_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a708_4 ( .OUT(na708_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a708_6 ( .RAM_O2(na708_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na708_2), .COMP_OUT(1'b0) );
// C_AND////      x28y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a709_1 ( .OUT(na709_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a709_6 ( .RAM_O1(na709_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na709_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y72     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a710_4 ( .OUT(na710_2), .IN1(1'b1), .IN2(na136_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a710_6 ( .RAM_O2(na710_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na710_2), .COMP_OUT(1'b0) );
// C_AND////      x37y72     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a711_1 ( .OUT(na711_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na135_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a711_6 ( .RAM_O1(na711_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na711_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y71     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a712_4 ( .OUT(na712_2), .IN1(na134_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a712_6 ( .RAM_O2(na712_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na712_2), .COMP_OUT(1'b0) );
// C_AND////      x37y71     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a713_1 ( .OUT(na713_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na133_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a713_6 ( .RAM_O1(na713_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na713_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y70     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a714_4 ( .OUT(na714_2), .IN1(1'b1), .IN2(na132_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a714_6 ( .RAM_O2(na714_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na714_2), .COMP_OUT(1'b0) );
// C_AND////      x37y70     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a715_1 ( .OUT(na715_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na131_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a715_6 ( .RAM_O1(na715_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na715_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y69     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a716_4 ( .OUT(na716_2), .IN1(1'b1), .IN2(1'b1), .IN3(na130_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a716_6 ( .RAM_O2(na716_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na716_2), .COMP_OUT(1'b0) );
// C_AND////      x37y69     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a717_1 ( .OUT(na717_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na129_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a717_6 ( .RAM_O1(na717_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na717_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y68     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a718_4 ( .OUT(na718_2), .IN1(1'b1), .IN2(na128_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a718_6 ( .RAM_O2(na718_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na718_2), .COMP_OUT(1'b0) );
// C_AND////      x37y68     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a719_1 ( .OUT(na719_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na127_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a719_6 ( .RAM_O1(na719_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na719_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y67     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a720_4 ( .OUT(na720_2), .IN1(1'b1), .IN2(na126_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a720_6 ( .RAM_O2(na720_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na720_2), .COMP_OUT(1'b0) );
// C_AND////      x37y67     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a721_1 ( .OUT(na721_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na125_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a721_6 ( .RAM_O1(na721_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na721_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y66     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a722_4 ( .OUT(na722_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na124_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a722_6 ( .RAM_O2(na722_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na722_2), .COMP_OUT(1'b0) );
// C_AND////      x37y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a723_1 ( .OUT(na723_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a723_6 ( .RAM_O1(na723_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na723_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a724_4 ( .OUT(na724_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a724_6 ( .RAM_O2(na724_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na724_2), .COMP_OUT(1'b0) );
// C_AND////      x37y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a725_1 ( .OUT(na725_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a725_6 ( .RAM_O1(na725_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na725_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y80     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a726_4 ( .OUT(na726_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a726_6 ( .RAM_O2(na726_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na726_2), .COMP_OUT(1'b0) );
// C_AND////      x30y80     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a727_1 ( .OUT(na727_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a727_6 ( .RAM_O1(na727_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na727_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y79     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a728_4 ( .OUT(na728_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a728_6 ( .RAM_O2(na728_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na728_2), .COMP_OUT(1'b0) );
// C_AND////      x30y79     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a729_1 ( .OUT(na729_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a729_6 ( .RAM_O1(na729_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na729_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y80     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a730_4 ( .OUT(na730_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a730_6 ( .RAM_O2(na730_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na730_2), .COMP_OUT(1'b0) );
// C_AND////      x32y80     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a731_1 ( .OUT(na731_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a731_6 ( .RAM_O1(na731_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na731_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y79     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a732_4 ( .OUT(na732_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a732_6 ( .RAM_O2(na732_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na732_2), .COMP_OUT(1'b0) );
// C_AND////      x32y79     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a733_1 ( .OUT(na733_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a733_6 ( .RAM_O1(na733_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na733_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y78     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a734_4 ( .OUT(na734_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a734_6 ( .RAM_O2(na734_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na734_2), .COMP_OUT(1'b0) );
// C_AND////      x32y78     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a735_1 ( .OUT(na735_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a735_6 ( .RAM_O1(na735_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na735_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y77     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a736_4 ( .OUT(na736_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a736_6 ( .RAM_O2(na736_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na736_2), .COMP_OUT(1'b0) );
// C_AND////      x32y77     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a737_1 ( .OUT(na737_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a737_6 ( .RAM_O1(na737_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na737_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y76     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a738_4 ( .OUT(na738_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a738_6 ( .RAM_O2(na738_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na738_2), .COMP_OUT(1'b0) );
// C_AND////      x32y76     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a739_1 ( .OUT(na739_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a739_6 ( .RAM_O1(na739_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na739_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y75     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a740_4 ( .OUT(na740_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a740_6 ( .RAM_O2(na740_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na740_2), .COMP_OUT(1'b0) );
// C_AND////      x32y75     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a741_1 ( .OUT(na741_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a741_6 ( .RAM_O1(na741_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na741_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y74     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a742_4 ( .OUT(na742_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a742_6 ( .RAM_O2(na742_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na742_2), .COMP_OUT(1'b0) );
// C_AND////      x32y74     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a743_1 ( .OUT(na743_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a743_6 ( .RAM_O1(na743_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na743_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y73     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a744_4 ( .OUT(na744_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a744_6 ( .RAM_O2(na744_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na744_2), .COMP_OUT(1'b0) );
// C_AND////      x32y73     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a745_1 ( .OUT(na745_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a745_6 ( .RAM_O1(na745_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na745_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a746_4 ( .OUT(na746_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a746_6 ( .RAM_O2(na746_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na746_2), .COMP_OUT(1'b0) );
// C_AND////      x30y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a747_1 ( .OUT(na747_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a747_6 ( .RAM_O1(na747_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na747_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a748_4 ( .OUT(na748_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a748_6 ( .RAM_O2(na748_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na748_2), .COMP_OUT(1'b0) );
// C_AND////      x30y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a749_1 ( .OUT(na749_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a749_6 ( .RAM_O1(na749_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na749_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a750_4 ( .OUT(na750_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a750_6 ( .RAM_O2(na750_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na750_2), .COMP_OUT(1'b0) );
// C_AND////      x32y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a751_1 ( .OUT(na751_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a751_6 ( .RAM_O1(na751_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na751_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a752_4 ( .OUT(na752_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a752_6 ( .RAM_O2(na752_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na752_2), .COMP_OUT(1'b0) );
// C_AND////      x32y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a753_1 ( .OUT(na753_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a753_6 ( .RAM_O1(na753_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na753_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y70     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a754_4 ( .OUT(na754_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a754_6 ( .RAM_O2(na754_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na754_2), .COMP_OUT(1'b0) );
// C_AND////      x32y70     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a755_1 ( .OUT(na755_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a755_6 ( .RAM_O1(na755_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na755_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y69     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a756_4 ( .OUT(na756_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a756_6 ( .RAM_O2(na756_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na756_2), .COMP_OUT(1'b0) );
// C_AND////      x32y69     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a757_1 ( .OUT(na757_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a757_6 ( .RAM_O1(na757_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na757_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y68     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a758_4 ( .OUT(na758_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a758_6 ( .RAM_O2(na758_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na758_2), .COMP_OUT(1'b0) );
// C_AND////      x32y68     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a759_1 ( .OUT(na759_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a759_6 ( .RAM_O1(na759_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na759_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y67     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a760_4 ( .OUT(na760_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a760_6 ( .RAM_O2(na760_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na760_2), .COMP_OUT(1'b0) );
// C_AND////      x32y67     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a761_1 ( .OUT(na761_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a761_6 ( .RAM_O1(na761_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na761_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y66     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a762_4 ( .OUT(na762_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a762_6 ( .RAM_O2(na762_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na762_2), .COMP_OUT(1'b0) );
// C_AND////      x32y66     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a763_1 ( .OUT(na763_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na390_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a763_6 ( .RAM_O1(na763_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na763_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y65     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a764_4 ( .OUT(na764_2), .IN1(1'b1), .IN2(na250_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a764_6 ( .RAM_O2(na764_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na764_2), .COMP_OUT(1'b0) );
// C_AND////      x32y65     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a765_1 ( .OUT(na765_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na403_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a765_6 ( .RAM_O1(na765_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na765_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y80     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a766_4 ( .OUT(na766_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a766_6 ( .RAM_O2(na766_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na766_2), .COMP_OUT(1'b0) );
// C_AND////      x29y80     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a767_1 ( .OUT(na767_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a767_6 ( .RAM_O1(na767_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na767_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y79     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a768_4 ( .OUT(na768_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a768_6 ( .RAM_O2(na768_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na768_2), .COMP_OUT(1'b0) );
// C_AND////      x29y79     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a769_1 ( .OUT(na769_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a769_6 ( .RAM_O1(na769_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na769_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y80     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a770_4 ( .OUT(na770_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a770_6 ( .RAM_O2(na770_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na770_2), .COMP_OUT(1'b0) );
// C_AND////      x31y80     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a771_1 ( .OUT(na771_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a771_6 ( .RAM_O1(na771_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na771_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y79     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a772_4 ( .OUT(na772_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a772_6 ( .RAM_O2(na772_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na772_2), .COMP_OUT(1'b0) );
// C_AND////      x31y79     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a773_1 ( .OUT(na773_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a773_6 ( .RAM_O1(na773_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na773_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y78     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a774_4 ( .OUT(na774_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a774_6 ( .RAM_O2(na774_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na774_2), .COMP_OUT(1'b0) );
// C_AND////      x31y78     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a775_1 ( .OUT(na775_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a775_6 ( .RAM_O1(na775_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na775_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y77     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a776_4 ( .OUT(na776_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a776_6 ( .RAM_O2(na776_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na776_2), .COMP_OUT(1'b0) );
// C_AND////      x31y77     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a777_1 ( .OUT(na777_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a777_6 ( .RAM_O1(na777_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na777_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y76     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a778_4 ( .OUT(na778_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a778_6 ( .RAM_O2(na778_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na778_2), .COMP_OUT(1'b0) );
// C_AND////      x31y76     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a779_1 ( .OUT(na779_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a779_6 ( .RAM_O1(na779_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na779_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y75     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a780_4 ( .OUT(na780_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a780_6 ( .RAM_O2(na780_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na780_2), .COMP_OUT(1'b0) );
// C_AND////      x31y75     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a781_1 ( .OUT(na781_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a781_6 ( .RAM_O1(na781_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na781_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y74     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a782_4 ( .OUT(na782_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a782_6 ( .RAM_O2(na782_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na782_2), .COMP_OUT(1'b0) );
// C_AND////      x31y74     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a783_1 ( .OUT(na783_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a783_6 ( .RAM_O1(na783_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na783_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y73     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a784_4 ( .OUT(na784_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a784_6 ( .RAM_O2(na784_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na784_2), .COMP_OUT(1'b0) );
// C_AND////      x31y73     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a785_1 ( .OUT(na785_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a785_6 ( .RAM_O1(na785_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na785_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a786_4 ( .OUT(na786_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a786_6 ( .RAM_O2(na786_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na786_2), .COMP_OUT(1'b0) );
// C_AND////      x29y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a787_1 ( .OUT(na787_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a787_6 ( .RAM_O1(na787_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na787_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a788_4 ( .OUT(na788_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a788_6 ( .RAM_O2(na788_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na788_2), .COMP_OUT(1'b0) );
// C_AND////      x29y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a789_1 ( .OUT(na789_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a789_6 ( .RAM_O1(na789_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na789_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a790_4 ( .OUT(na790_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a790_6 ( .RAM_O2(na790_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na790_2), .COMP_OUT(1'b0) );
// C_AND////      x31y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a791_1 ( .OUT(na791_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a791_6 ( .RAM_O1(na791_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na791_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a792_4 ( .OUT(na792_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a792_6 ( .RAM_O2(na792_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na792_2), .COMP_OUT(1'b0) );
// C_AND////      x31y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a793_1 ( .OUT(na793_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a793_6 ( .RAM_O1(na793_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na793_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y70     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a794_4 ( .OUT(na794_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a794_6 ( .RAM_O2(na794_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na794_2), .COMP_OUT(1'b0) );
// C_AND////      x31y70     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a795_1 ( .OUT(na795_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a795_6 ( .RAM_O1(na795_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na795_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y69     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a796_4 ( .OUT(na796_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a796_6 ( .RAM_O2(na796_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na796_2), .COMP_OUT(1'b0) );
// C_AND////      x31y69     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a797_1 ( .OUT(na797_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a797_6 ( .RAM_O1(na797_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na797_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y68     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a798_4 ( .OUT(na798_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a798_6 ( .RAM_O2(na798_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na798_2), .COMP_OUT(1'b0) );
// C_AND////      x31y68     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a799_1 ( .OUT(na799_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a799_6 ( .RAM_O1(na799_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na799_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y67     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a800_4 ( .OUT(na800_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a800_6 ( .RAM_O2(na800_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na800_2), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x34y66     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a801_2 ( .OUT(na801_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na400_118), .CP_O(1'b0) );
// C_////RAM_I2      x34y65     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a802_5 ( .OUT(na802_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na400_119), .CP_O(1'b0) );
// C_/RAM_I1///      x34y65     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a803_2 ( .OUT(na803_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na400_120), .CP_O(1'b0) );
// C_AND////      x35y17     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a804_1 ( .OUT(na804_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na392_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a804_6 ( .RAM_O1(na804_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na804_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x27y17     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a805_4 ( .OUT(na805_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na147_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a805_6 ( .RAM_O2(na805_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na805_2), .COMP_OUT(1'b0) );
// C_///AND/      x28y24     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a806_4 ( .OUT(na806_2), .IN1(1'b1), .IN2(na97_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a806_6 ( .RAM_O2(na806_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na806_2), .COMP_OUT(1'b0) );
// C_AND////      x28y24     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a807_1 ( .OUT(na807_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na97_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a807_6 ( .RAM_O1(na807_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na807_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y23     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a808_4 ( .OUT(na808_2), .IN1(1'b1), .IN2(na99_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a808_6 ( .RAM_O2(na808_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na808_2), .COMP_OUT(1'b0) );
// C_AND////      x28y23     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a809_1 ( .OUT(na809_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na99_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a809_6 ( .RAM_O1(na809_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na809_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y22     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a810_4 ( .OUT(na810_2), .IN1(na84_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a810_6 ( .RAM_O2(na810_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na810_2), .COMP_OUT(1'b0) );
// C_AND////      x28y22     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a811_1 ( .OUT(na811_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na84_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a811_6 ( .RAM_O1(na811_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na811_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y21     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a812_4 ( .OUT(na812_2), .IN1(1'b1), .IN2(na102_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a812_6 ( .RAM_O2(na812_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na812_2), .COMP_OUT(1'b0) );
// C_AND////      x28y21     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a813_1 ( .OUT(na813_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na102_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a813_6 ( .RAM_O1(na813_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na813_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y20     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a814_4 ( .OUT(na814_2), .IN1(na117_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a814_6 ( .RAM_O2(na814_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na814_2), .COMP_OUT(1'b0) );
// C_AND////      x28y20     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a815_1 ( .OUT(na815_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na117_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a815_6 ( .RAM_O1(na815_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na815_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y19     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a816_4 ( .OUT(na816_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a816_6 ( .RAM_O2(na816_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na816_2), .COMP_OUT(1'b0) );
// C_AND////      x28y19     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a817_1 ( .OUT(na817_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na8_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a817_6 ( .RAM_O1(na817_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na817_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y18     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a818_4 ( .OUT(na818_2), .IN1(1'b1), .IN2(1'b1), .IN3(na15_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a818_6 ( .RAM_O2(na818_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na818_2), .COMP_OUT(1'b0) );
// C_AND////      x28y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a819_1 ( .OUT(na819_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a819_6 ( .RAM_O1(na819_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na819_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a820_4 ( .OUT(na820_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a820_6 ( .RAM_O2(na820_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na820_2), .COMP_OUT(1'b0) );
// C_AND////      x28y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a821_1 ( .OUT(na821_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a821_6 ( .RAM_O1(na821_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na821_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y24     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a822_4 ( .OUT(na822_2), .IN1(1'b1), .IN2(na136_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a822_6 ( .RAM_O2(na822_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na822_2), .COMP_OUT(1'b0) );
// C_AND////      x37y24     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a823_1 ( .OUT(na823_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na135_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a823_6 ( .RAM_O1(na823_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na823_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y23     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a824_4 ( .OUT(na824_2), .IN1(na134_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a824_6 ( .RAM_O2(na824_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na824_2), .COMP_OUT(1'b0) );
// C_AND////      x37y23     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a825_1 ( .OUT(na825_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na133_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a825_6 ( .RAM_O1(na825_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na825_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y22     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a826_4 ( .OUT(na826_2), .IN1(1'b1), .IN2(na132_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a826_6 ( .RAM_O2(na826_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na826_2), .COMP_OUT(1'b0) );
// C_AND////      x37y22     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a827_1 ( .OUT(na827_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na131_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a827_6 ( .RAM_O1(na827_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na827_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y21     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a828_4 ( .OUT(na828_2), .IN1(1'b1), .IN2(1'b1), .IN3(na130_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a828_6 ( .RAM_O2(na828_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na828_2), .COMP_OUT(1'b0) );
// C_AND////      x37y21     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a829_1 ( .OUT(na829_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na129_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a829_6 ( .RAM_O1(na829_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na829_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y20     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a830_4 ( .OUT(na830_2), .IN1(1'b1), .IN2(na128_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a830_6 ( .RAM_O2(na830_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na830_2), .COMP_OUT(1'b0) );
// C_AND////      x37y20     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a831_1 ( .OUT(na831_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na127_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a831_6 ( .RAM_O1(na831_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na831_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y19     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a832_4 ( .OUT(na832_2), .IN1(1'b1), .IN2(na126_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a832_6 ( .RAM_O2(na832_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na832_2), .COMP_OUT(1'b0) );
// C_AND////      x37y19     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a833_1 ( .OUT(na833_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na125_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a833_6 ( .RAM_O1(na833_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na833_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y18     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a834_4 ( .OUT(na834_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na124_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a834_6 ( .RAM_O2(na834_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na834_2), .COMP_OUT(1'b0) );
// C_AND////      x37y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a835_1 ( .OUT(na835_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a835_6 ( .RAM_O1(na835_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na835_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a836_4 ( .OUT(na836_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a836_6 ( .RAM_O2(na836_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na836_2), .COMP_OUT(1'b0) );
// C_AND////      x37y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a837_1 ( .OUT(na837_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a837_6 ( .RAM_O1(na837_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na837_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y32     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a838_4 ( .OUT(na838_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a838_6 ( .RAM_O2(na838_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na838_2), .COMP_OUT(1'b0) );
// C_AND////      x30y32     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a839_1 ( .OUT(na839_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a839_6 ( .RAM_O1(na839_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na839_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y31     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a840_4 ( .OUT(na840_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a840_6 ( .RAM_O2(na840_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na840_2), .COMP_OUT(1'b0) );
// C_AND////      x30y31     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a841_1 ( .OUT(na841_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a841_6 ( .RAM_O1(na841_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na841_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y32     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a842_4 ( .OUT(na842_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a842_6 ( .RAM_O2(na842_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na842_2), .COMP_OUT(1'b0) );
// C_AND////      x32y32     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a843_1 ( .OUT(na843_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a843_6 ( .RAM_O1(na843_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na843_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y31     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a844_4 ( .OUT(na844_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a844_6 ( .RAM_O2(na844_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na844_2), .COMP_OUT(1'b0) );
// C_AND////      x32y31     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a845_1 ( .OUT(na845_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a845_6 ( .RAM_O1(na845_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na845_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y30     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a846_4 ( .OUT(na846_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a846_6 ( .RAM_O2(na846_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na846_2), .COMP_OUT(1'b0) );
// C_AND////      x32y30     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a847_1 ( .OUT(na847_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a847_6 ( .RAM_O1(na847_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na847_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y29     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a848_4 ( .OUT(na848_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a848_6 ( .RAM_O2(na848_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na848_2), .COMP_OUT(1'b0) );
// C_AND////      x32y29     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a849_1 ( .OUT(na849_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a849_6 ( .RAM_O1(na849_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na849_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y28     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a850_4 ( .OUT(na850_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a850_6 ( .RAM_O2(na850_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na850_2), .COMP_OUT(1'b0) );
// C_AND////      x32y28     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a851_1 ( .OUT(na851_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a851_6 ( .RAM_O1(na851_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na851_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y27     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a852_4 ( .OUT(na852_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a852_6 ( .RAM_O2(na852_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na852_2), .COMP_OUT(1'b0) );
// C_AND////      x32y27     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a853_1 ( .OUT(na853_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a853_6 ( .RAM_O1(na853_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na853_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y26     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a854_4 ( .OUT(na854_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a854_6 ( .RAM_O2(na854_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na854_2), .COMP_OUT(1'b0) );
// C_AND////      x32y26     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a855_1 ( .OUT(na855_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a855_6 ( .RAM_O1(na855_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na855_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y25     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a856_4 ( .OUT(na856_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a856_6 ( .RAM_O2(na856_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na856_2), .COMP_OUT(1'b0) );
// C_AND////      x32y25     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a857_1 ( .OUT(na857_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a857_6 ( .RAM_O1(na857_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na857_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y24     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a858_4 ( .OUT(na858_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a858_6 ( .RAM_O2(na858_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na858_2), .COMP_OUT(1'b0) );
// C_AND////      x30y24     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a859_1 ( .OUT(na859_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a859_6 ( .RAM_O1(na859_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na859_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y23     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a860_4 ( .OUT(na860_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a860_6 ( .RAM_O2(na860_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na860_2), .COMP_OUT(1'b0) );
// C_AND////      x30y23     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a861_1 ( .OUT(na861_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a861_6 ( .RAM_O1(na861_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na861_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y24     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a862_4 ( .OUT(na862_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a862_6 ( .RAM_O2(na862_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na862_2), .COMP_OUT(1'b0) );
// C_AND////      x32y24     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a863_1 ( .OUT(na863_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a863_6 ( .RAM_O1(na863_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na863_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y23     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a864_4 ( .OUT(na864_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a864_6 ( .RAM_O2(na864_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na864_2), .COMP_OUT(1'b0) );
// C_AND////      x32y23     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a865_1 ( .OUT(na865_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a865_6 ( .RAM_O1(na865_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na865_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y22     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a866_4 ( .OUT(na866_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a866_6 ( .RAM_O2(na866_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na866_2), .COMP_OUT(1'b0) );
// C_AND////      x32y22     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a867_1 ( .OUT(na867_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a867_6 ( .RAM_O1(na867_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na867_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y21     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a868_4 ( .OUT(na868_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a868_6 ( .RAM_O2(na868_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na868_2), .COMP_OUT(1'b0) );
// C_AND////      x32y21     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a869_1 ( .OUT(na869_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a869_6 ( .RAM_O1(na869_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na869_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y20     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a870_4 ( .OUT(na870_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a870_6 ( .RAM_O2(na870_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na870_2), .COMP_OUT(1'b0) );
// C_AND////      x32y20     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a871_1 ( .OUT(na871_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a871_6 ( .RAM_O1(na871_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na871_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y19     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a872_4 ( .OUT(na872_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a872_6 ( .RAM_O2(na872_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na872_2), .COMP_OUT(1'b0) );
// C_AND////      x32y19     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a873_1 ( .OUT(na873_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a873_6 ( .RAM_O1(na873_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na873_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y18     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a874_4 ( .OUT(na874_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a874_6 ( .RAM_O2(na874_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na874_2), .COMP_OUT(1'b0) );
// C_AND////      x32y18     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a875_1 ( .OUT(na875_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na390_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a875_6 ( .RAM_O1(na875_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na875_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y17     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a876_4 ( .OUT(na876_2), .IN1(1'b1), .IN2(na250_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a876_6 ( .RAM_O2(na876_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na876_2), .COMP_OUT(1'b0) );
// C_AND////      x32y17     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a877_1 ( .OUT(na877_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na403_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a877_6 ( .RAM_O1(na877_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na877_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y32     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a878_4 ( .OUT(na878_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a878_6 ( .RAM_O2(na878_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na878_2), .COMP_OUT(1'b0) );
// C_AND////      x29y32     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a879_1 ( .OUT(na879_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a879_6 ( .RAM_O1(na879_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na879_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y31     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a880_4 ( .OUT(na880_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a880_6 ( .RAM_O2(na880_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na880_2), .COMP_OUT(1'b0) );
// C_AND////      x29y31     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a881_1 ( .OUT(na881_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a881_6 ( .RAM_O1(na881_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na881_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y32     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a882_4 ( .OUT(na882_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a882_6 ( .RAM_O2(na882_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na882_2), .COMP_OUT(1'b0) );
// C_AND////      x31y32     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a883_1 ( .OUT(na883_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a883_6 ( .RAM_O1(na883_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na883_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y31     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a884_4 ( .OUT(na884_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a884_6 ( .RAM_O2(na884_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na884_2), .COMP_OUT(1'b0) );
// C_AND////      x31y31     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a885_1 ( .OUT(na885_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a885_6 ( .RAM_O1(na885_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na885_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y30     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a886_4 ( .OUT(na886_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a886_6 ( .RAM_O2(na886_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na886_2), .COMP_OUT(1'b0) );
// C_AND////      x31y30     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a887_1 ( .OUT(na887_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a887_6 ( .RAM_O1(na887_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na887_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y29     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a888_4 ( .OUT(na888_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a888_6 ( .RAM_O2(na888_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na888_2), .COMP_OUT(1'b0) );
// C_AND////      x31y29     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a889_1 ( .OUT(na889_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a889_6 ( .RAM_O1(na889_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na889_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y28     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a890_4 ( .OUT(na890_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a890_6 ( .RAM_O2(na890_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na890_2), .COMP_OUT(1'b0) );
// C_AND////      x31y28     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a891_1 ( .OUT(na891_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a891_6 ( .RAM_O1(na891_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na891_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y27     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a892_4 ( .OUT(na892_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a892_6 ( .RAM_O2(na892_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na892_2), .COMP_OUT(1'b0) );
// C_AND////      x31y27     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a893_1 ( .OUT(na893_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a893_6 ( .RAM_O1(na893_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na893_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y26     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a894_4 ( .OUT(na894_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a894_6 ( .RAM_O2(na894_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na894_2), .COMP_OUT(1'b0) );
// C_AND////      x31y26     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a895_1 ( .OUT(na895_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a895_6 ( .RAM_O1(na895_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na895_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y25     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a896_4 ( .OUT(na896_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a896_6 ( .RAM_O2(na896_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na896_2), .COMP_OUT(1'b0) );
// C_AND////      x31y25     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a897_1 ( .OUT(na897_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a897_6 ( .RAM_O1(na897_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na897_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y24     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a898_4 ( .OUT(na898_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a898_6 ( .RAM_O2(na898_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na898_2), .COMP_OUT(1'b0) );
// C_AND////      x29y24     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a899_1 ( .OUT(na899_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a899_6 ( .RAM_O1(na899_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na899_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y23     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a900_4 ( .OUT(na900_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a900_6 ( .RAM_O2(na900_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na900_2), .COMP_OUT(1'b0) );
// C_AND////      x29y23     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a901_1 ( .OUT(na901_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a901_6 ( .RAM_O1(na901_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na901_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y24     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a902_4 ( .OUT(na902_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a902_6 ( .RAM_O2(na902_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na902_2), .COMP_OUT(1'b0) );
// C_AND////      x31y24     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a903_1 ( .OUT(na903_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a903_6 ( .RAM_O1(na903_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na903_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y23     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a904_4 ( .OUT(na904_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a904_6 ( .RAM_O2(na904_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na904_2), .COMP_OUT(1'b0) );
// C_AND////      x31y23     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a905_1 ( .OUT(na905_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a905_6 ( .RAM_O1(na905_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na905_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y22     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a906_4 ( .OUT(na906_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a906_6 ( .RAM_O2(na906_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na906_2), .COMP_OUT(1'b0) );
// C_AND////      x31y22     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a907_1 ( .OUT(na907_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a907_6 ( .RAM_O1(na907_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na907_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y21     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a908_4 ( .OUT(na908_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a908_6 ( .RAM_O2(na908_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na908_2), .COMP_OUT(1'b0) );
// C_AND////      x31y21     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a909_1 ( .OUT(na909_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a909_6 ( .RAM_O1(na909_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na909_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y20     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a910_4 ( .OUT(na910_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a910_6 ( .RAM_O2(na910_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na910_2), .COMP_OUT(1'b0) );
// C_AND////      x31y20     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a911_1 ( .OUT(na911_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a911_6 ( .RAM_O1(na911_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na911_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y19     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a912_4 ( .OUT(na912_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a912_6 ( .RAM_O2(na912_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na912_2), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x34y18     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a913_2 ( .OUT(na913_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na401_118), .CP_O(1'b0) );
// C_////RAM_I2      x34y17     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a914_5 ( .OUT(na914_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na401_119), .CP_O(1'b0) );
// C_/RAM_I1///      x34y17     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a915_2 ( .OUT(na915_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na401_120), .CP_O(1'b0) );
// C_////Bridge      x44y42     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a916_5 ( .OUT(na916_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y41     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a917_5 ( .OUT(na917_2), .IN1(1'b0), .IN2(na1_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y45     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a918_5 ( .OUT(na918_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y44     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a919_5 ( .OUT(na919_2), .IN1(1'b0), .IN2(1'b0), .IN3(na4_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y44     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a920_5 ( .OUT(na920_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na6_1) );
// C_////Bridge      x47y44     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a921_5 ( .OUT(na921_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na6_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y43     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a922_5 ( .OUT(na922_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y39     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a923_5 ( .OUT(na923_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na7_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y54     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a924_5 ( .OUT(na924_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na13_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y51     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a925_5 ( .OUT(na925_2), .IN1(1'b0), .IN2(na14_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y40     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a926_5 ( .OUT(na926_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na17_1) );
// C_////Bridge      x47y42     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a927_5 ( .OUT(na927_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na17_2) );
// C_////Bridge      x36y39     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a928_5 ( .OUT(na928_2), .IN1(na25_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y42     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a929_5 ( .OUT(na929_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na27_2), .IN8(1'b0) );
// C_////Bridge      x36y42     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a930_5 ( .OUT(na930_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na31_2), .IN8(1'b0) );
// C_////Bridge      x39y43     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a931_5 ( .OUT(na931_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na87_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y37     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a932_5 ( .OUT(na932_2), .IN1(1'b0), .IN2(1'b0), .IN3(na91_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y51     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a933_5 ( .OUT(na933_2), .IN1(1'b0), .IN2(1'b0), .IN3(na91_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y37     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a934_5 ( .OUT(na934_2), .IN1(1'b0), .IN2(1'b0), .IN3(na93_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y42     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a935_5 ( .OUT(na935_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na112_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a936_5 ( .OUT(na936_2), .IN1(1'b0), .IN2(1'b0), .IN3(na113_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y49     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a937_5 ( .OUT(na937_2), .IN1(na137_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y40     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a938_5 ( .OUT(na938_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na140_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y39     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a939_5 ( .OUT(na939_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na156_2), .IN8(1'b0) );
// C_////Bridge      x42y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a940_5 ( .OUT(na940_2), .IN1(1'b0), .IN2(1'b0), .IN3(na190_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y48     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a941_5 ( .OUT(na941_2), .IN1(1'b0), .IN2(1'b0), .IN3(na190_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y46     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a942_5 ( .OUT(na942_2), .IN1(1'b0), .IN2(1'b0), .IN3(na196_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y46     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a943_5 ( .OUT(na943_2), .IN1(1'b0), .IN2(1'b0), .IN3(na196_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y44     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a944_5 ( .OUT(na944_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na200_1), .IN8(1'b0) );
// C_////Bridge      x36y44     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a945_5 ( .OUT(na945_2), .IN1(1'b0), .IN2(1'b0), .IN3(na200_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y47     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a946_5 ( .OUT(na946_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na207_1) );
// C_////Bridge      x40y39     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a947_5 ( .OUT(na947_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na207_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y39     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a948_5 ( .OUT(na948_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na209_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y41     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a949_5 ( .OUT(na949_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na209_2) );
// C_////Bridge      x42y43     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a950_5 ( .OUT(na950_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na213_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y47     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a951_5 ( .OUT(na951_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na213_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y45     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a952_5 ( .OUT(na952_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na217_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y45     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a953_5 ( .OUT(na953_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na217_2) );
// C_////Bridge      x42y53     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a954_5 ( .OUT(na954_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na577_1) );
// C_////Bridge      x38y32     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a955_5 ( .OUT(na955_2), .IN1(1'b0), .IN2(1'b0), .IN3(na690_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y34     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a956_5 ( .OUT(na956_2), .IN1(1'b0), .IN2(1'b0), .IN3(na691_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y52     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a957_5 ( .OUT(na957_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na802_2), .IN8(1'b0) );
// C_////Bridge      x34y46     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a958_5 ( .OUT(na958_2), .IN1(1'b0), .IN2(1'b0), .IN3(na803_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y35     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a959_5 ( .OUT(na959_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na913_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
endmodule
