//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 July 2024)
//  Compile Time: 2024-07-19 13:57:40
//  Program Run:  2024-08-31 21:45:56
//  Program Call: /home/user/FPGA/Boards/GateMate/cc-toolchain-linux//bin/p_r/p_r -i net/top_synth.v -o top -ccf /home/user/openCologne/10.Bonus--4--I2C-Master/3.build/../1.hw/constraints/top.ccf -cCP 
//  File Type:    Verilog

// Gatecount:    232
module top (areset_n , clk_10MHz ,
       led ,
       i2c_scl , i2c_sda 
) ;

input  areset_n;
input  clk_10MHz;

output led;

inout  i2c_scl;
inout  i2c_sda;


wire led;
wire na1_1;
wire na2_1;
wire na2_2;
wire na4_1;
wire na4_1_i;
wire na4_2;
wire na4_2_i;
wire na5_1;
wire na5_1_i;
wire na5_2;
wire na5_2_i;
wire na8_1;
wire na8_1_i;
wire na8_2;
wire na8_2_i;
wire na9_2;
wire na9_2_i;
wire na10_1;
wire na10_1_i;
wire na12_1;
wire na13_1;
wire na14_2;
wire na15_1;
wire na15_1_i;
wire na16_1;
wire na19_1;
wire na20_1;
wire na21_1;
wire na21_2;
wire na22_1;
wire na22_2;
wire na23_2;
wire na23_2_i;
wire na24_1;
wire na24_1_i;
wire na26_1;
wire na27_1;
wire na28_1;
wire na28_1_i;
wire na29_2;
wire na29_2_i;
wire na31_1;
wire na31_1_i;
wire na32_1;
wire na32_1_i;
wire na32_2;
wire na32_2_i;
wire na33_2;
wire na33_2_i;
wire na35_1;
wire na36_1;
wire na37_2;
wire na38_2;
wire na39_1;
wire na40_2;
wire na42_1;
wire na43_1;
wire na44_1;
wire na44_2;
wire na45_2;
wire na46_2;
wire na47_1;
wire na48_1;
wire na49_1;
wire na51_2;
wire na52_1;
wire na53_2;
wire na54_1;
wire na55_1;
wire na56_2;
wire na57_1;
wire na58_1;
wire na59_1;
wire na60_2;
wire na61_2;
wire na61_2_i;
wire na62_1;
wire na62_1_i;
wire na63_1;
wire na65_1;
wire na66_1;
wire na66_2;
wire na67_1;
wire na70_1;
wire na71_1;
wire na71_1_i;
wire na72_1;
wire na72_1_i;
wire na74_2;
wire na74_2_i;
wire na75_1;
wire na77_1;
wire na77_1_i;
wire na78_2;
wire na78_2_i;
wire na79_2;
wire na80_1;
wire na81_1;
wire na83_1;
wire na84_2;
wire na85_1;
wire na88_1;
wire na89_1;
wire na90_1;
wire na91_1;
wire na92_2;
wire na93_2;
wire na94_1;
wire i2c_scl;
wire i2c_sda;
wire na102_1;
wire na103_1;
wire na104_1;
wire na105_1;
wire na106_1;
wire na107_1;
wire na108_1;
wire na110_4;
wire na112_4;
wire na114_4;
wire na116_1;
wire na116_4;
wire na117_1;
wire na117_2;
wire na117_4;
wire na119_1;
wire na119_2;
wire na119_4;
wire na121_1;
wire na121_2;
wire na123_1;
wire na123_4;
wire na125_1;
wire na125_1_i;
wire na125_2;
wire na125_4;
wire na127_1;
wire na127_1_i;
wire na127_2;
wire na127_4;
wire na129_1;
wire na129_1_i;
wire na129_2;
wire na129_4;
wire na131_1;
wire na131_1_i;
wire na131_2;
wire na131_4;
wire na133_1;
wire na133_1_i;
wire na133_2;
wire na133_4;
wire na134_1;
wire na134_1_i;
wire na134_2;
wire na134_4;
wire na136_1;
wire na136_1_i;
wire na136_2;
wire na136_4;
wire na138_1;
wire na138_1_i;
wire na140_1;
wire na140_1_i;
wire na140_2;
wire na140_4;
wire na142_1;
wire na142_1_i;
wire na142_2;
wire na142_4;
wire na144_1;
wire na144_1_i;
wire na144_2;
wire na144_4;
wire na146_1;
wire na146_1_i;
wire na146_2;
wire na146_4;
wire na147_1;
wire na147_4;
wire na148_1;
wire na148_1_i;
wire na148_2;
wire na148_4;
wire na150_1;
wire na150_1_i;
wire na150_2;
wire na150_4;
wire na152_1;
wire na152_1_i;
wire na152_2;
wire na154_1;
wire na154_4;
wire na155_1;
wire na155_2;
wire na155_4;
wire na157_1;
wire na158_1;
wire na158_4;
wire na159_1;
wire na159_2;
wire na159_4;
wire na161_1;
wire na163_1;
wire na165_1;
wire na165_1_i;
wire na165_2;
wire na165_2_i;
wire na167_2;
wire na167_2_i;
wire na169_1;
wire na169_1_i;
wire na171_2;
wire na171_2_i;
wire na173_1;
wire na173_1_i;
wire na175_2;
wire na175_2_i;
wire na177_2;
wire na177_2_i;
wire na179_1;
wire na179_1_i;
wire na181_2;
wire na181_2_i;
wire na183_1;
wire na183_1_i;
wire na185_1;
wire na185_1_i;
wire na214_2;
wire na214_2_i;
wire na218_1;
wire na218_1_i;
wire na218_2;
wire na218_2_i;
wire na220_1;
wire na220_1_i;
wire na222_1;
wire na223_1;
wire na224_1;
wire na225_1;
wire na226_1;
wire na227_1;
wire na228_1;
wire na229_1;
wire na230_1;
wire na231_1;
wire na232_1;
wire na233_1;
wire na234_1;
wire na235_1;
wire na236_1;
wire na237_1;
wire na238_1;
wire na239_1;
wire na240_1;
wire na241_1;
wire na242_1;
wire na243_1;
wire na244_1;
wire na245_1;
wire na248_1;
wire na249_1;
wire na249_2;
wire na250_2;
wire na250_2_i;
wire na252_2;
wire na253_1;
wire na254_1;
wire na256_1;
wire na258_2;
wire na259_2;
wire na260_1;
wire na260_4;
wire na262_2;
wire na266_2;
wire na272_1;
wire na273_1;
wire na275_1;
wire na276_1;
wire na277_1;
wire na278_1;
wire na280_1;
wire na282_1;
wire na283_1;
wire na284_1;
wire na284_2;
wire na286_1;
wire na288_2;
wire na289_1;
wire na290_2;
wire na292_2;
wire na294_2;
wire na295_2;
wire na296_2;
wire na297_2;
wire na298_2;
wire na299_2;
wire na300_2;
wire na301_2;
wire na302_2;
wire na303_2;
wire na304_2;
wire na305_2;
wire na306_2;
wire na307_2;
wire na308_2;
wire na309_2;
wire na310_2;
wire na311_2;
wire na312_2;
wire na313_2;
wire na314_2;
wire na315_2;
wire na316_2;
wire na317_2;
wire na318_2;
wire na319_2;
wire na320_2;
wire na321_2;
wire na322_2;
wire na323_2;
wire na324_2;
wire na325_2;
wire na326_2;
wire na327_2;
wire na328_2;
wire na329_2;
wire na330_2;
wire na331_2;
wire na332_2;
wire na333_2;
wire na334_2;
wire na335_2;
wire na336_2;
wire na337_2;
wire na338_2;
wire na339_2;
wire na340_2;
wire na341_2;
wire na342_2;
wire na343_2;
wire na344_2;
wire na345_2;
wire na346_2;
wire na347_2;
wire areset_n;
wire na296_10;
wire na297_10;
wire na298_10;
wire na299_10;
wire na300_10;
wire clk_10MHz;

CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a1 ( .PCLK0(na1_1), .PCLK1(_d0), .PCLK2(_d1), .PCLK3(_d2), .CLK0(na245_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0), .SER_CLK(1'b0),
                 .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_AND////D      x30y120     80'h00_EE18_00_0000_0888_5248
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2_1 ( .OUT(na2_1), .IN1(na8_1), .IN2(na4_1), .IN3(~na5_1), .IN4(na9_2), .IN5(na8_2), .IN6(~na4_2), .IN7(~na5_2), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2_5 ( .OUT(na2_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2_1) );
// C_AND/D//AND/D      x29y122     80'h00_EE00_80_0000_0C88_3A3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4_1 ( .OUT(na4_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na117_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na2_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4_2 ( .OUT(na4_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4_4 ( .OUT(na4_2_i), .IN1(1'b1), .IN2(na119_2), .IN3(1'b1), .IN4(~na2_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4_5 ( .OUT(na4_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4_2_i) );
// C_AND/D//AND/D      x30y123     80'h00_EE00_80_0000_0C88_3A3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5_1 ( .OUT(na5_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na117_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na2_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5_2 ( .OUT(na5_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5_4 ( .OUT(na5_2_i), .IN1(1'b1), .IN2(na119_1), .IN3(1'b1), .IN4(~na2_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a5_5 ( .OUT(na5_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5_2_i) );
// C_AND/D//AND/D      x31y117     80'h00_EE00_80_0000_0C88_3A35
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na121_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na2_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a8_2 ( .OUT(na8_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na8_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8_4 ( .OUT(na8_2_i), .IN1(~na8_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a8_5 ( .OUT(na8_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na8_2_i) );
// C_///AND/D      x32y126     80'h00_EE00_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9_4 ( .OUT(na9_2_i), .IN1(na121_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a9_5 ( .OUT(na9_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na9_2_i) );
// C_AND*/DST///      x43y122     80'h20_BA00_00_0000_0388_C5FF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a10_1 ( .OUT(na10_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na66_2), .IN6(1'b1), .IN7(1'b1), .IN8(na13_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0100_0000)) 
           _a10_2 ( .OUT(na10_1), .CLK(na163_1), .EN(na93_2), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na10_1_i) );
// C_AND////      x36y116     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na28_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na29_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x38y116     80'h00_0018_00_0040_0C16_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1), .IN1(1'b1), .IN2(na330_2), .IN3(na74_2), .IN4(1'b0), .IN5(na28_1), .IN6(1'b1), .IN7(1'b1), .IN8(na29_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x36y112     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a14_4 ( .OUT(na14_2), .IN1(1'b1), .IN2(na32_2), .IN3(na250_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/DST///      x42y114     80'h20_BA00_00_0000_0788_75A3
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a15_1 ( .OUT(na15_1_i), .IN1(1'b0), .IN2(~na19_1), .IN3(na16_1), .IN4(1'b0), .IN5(~na20_1), .IN6(1'b0), .IN7(~na231_1),
                    .IN8(~na21_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0100_0000)) 
           _a15_2 ( .OUT(na15_1), .CLK(na163_1), .EN(na108_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na15_1_i) );
// C_MX2b////      x42y117     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a16_1 ( .OUT(na16_1), .IN1(1'b1), .IN2(~na249_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na226_1), .IN6(~na249_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x37y116     80'h00_0018_00_0040_0C62_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a19_1 ( .OUT(na19_1), .IN1(1'b0), .IN2(~na24_1), .IN3(1'b1), .IN4(1'b0), .IN5(~na28_1), .IN6(1'b1), .IN7(1'b1), .IN8(na29_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x33y115     80'h00_0018_00_0000_0C88_A8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a20_1 ( .OUT(na20_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na28_1), .IN6(na24_1), .IN7(na61_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x40y116     80'h00_EA18_00_0000_0888_F1CF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a21_1 ( .OUT(na21_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na29_2), .IN5(~na28_1), .IN6(~na24_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a21_5 ( .OUT(na21_2), .CLK(na163_1), .EN(na63_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na21_1) );
// C_MX4a////D      x36y113     80'h00_EA18_00_0040_0C62_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1), .IN1(1'b0), .IN2(~na24_1), .IN3(1'b1), .IN4(1'b0), .IN5(na28_1), .IN6(1'b1), .IN7(1'b1), .IN8(na29_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a22_5 ( .OUT(na22_2), .CLK(na163_1), .EN(na63_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na22_1) );
// C_///ORAND*/D      x41y118     80'h00_EA00_80_0000_0C07_FFA7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a23_4 ( .OUT(na23_2_i), .IN1(~na310_2), .IN2(~na24_1), .IN3(na22_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a23_5 ( .OUT(na23_2), .CLK(na163_1), .EN(na63_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na23_2_i) );
// C_ORAND*/D///      x35y120     80'h00_EA00_00_0000_0388_E5FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a24_1 ( .OUT(na24_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na66_2), .IN6(1'b0), .IN7(na27_1), .IN8(na252_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a24_2 ( .OUT(na24_1), .CLK(na163_1), .EN(na90_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na24_1_i) );
// C_AND////      x40y113     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a26_1 ( .OUT(na26_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na28_1), .IN6(~na62_1), .IN7(na307_2), .IN8(~na29_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x40y121     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na28_1), .IN6(1'b1), .IN7(1'b1), .IN8(na29_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x37y117     80'h00_EA00_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a28_1 ( .OUT(na28_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na304_2), .IN6(~na253_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a28_2 ( .OUT(na28_1), .CLK(na163_1), .EN(na90_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na28_1_i) );
// C_///OR/D      x38y118     80'h00_EA00_80_0000_0C0E_FFAC
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a29_4 ( .OUT(na29_2_i), .IN1(1'b0), .IN2(na254_1), .IN3(na26_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a29_5 ( .OUT(na29_2), .CLK(na163_1), .EN(na90_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na29_2_i) );
// C_AND/D///      x44y119     80'h00_EA00_00_0000_0C88_85FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a31_1 ( .OUT(na31_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na78_2), .IN6(1'b1), .IN7(na22_1), .IN8(na159_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a31_2 ( .OUT(na31_1), .CLK(na163_1), .EN(na81_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na31_1_i) );
// C_AND/D//AND/D      x37y118     80'h00_EA00_80_0000_0C88_85A1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a32_1 ( .OUT(na32_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na78_2), .IN6(1'b1), .IN7(na22_1), .IN8(na159_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a32_2 ( .OUT(na32_1), .CLK(na163_1), .EN(na81_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na32_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a32_4 ( .OUT(na32_2_i), .IN1(~na78_2), .IN2(~na32_2), .IN3(na22_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a32_5 ( .OUT(na32_2), .CLK(na163_1), .EN(na81_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na32_2_i) );
// C_///ORAND*/D      x36y118     80'h00_EA00_80_0000_0C07_FFD7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a33_4 ( .OUT(na33_2_i), .IN1(~na303_2), .IN2(~na24_1), .IN3(~na22_1), .IN4(na256_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a33_5 ( .OUT(na33_2), .CLK(na163_1), .EN(na81_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na33_2_i) );
// C_AND////      x36y122     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a35_1 ( .OUT(na35_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na214_2), .IN6(~na148_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x36y120     80'h00_0018_00_0000_0C66_0600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na214_2), .IN6(na148_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x35y118     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a37_4 ( .OUT(na37_2), .IN1(1'b1), .IN2(~na345_2), .IN3(1'b1), .IN4(na36_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x35y119     80'h00_0060_00_0000_0C08_FFE3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a38_4 ( .OUT(na38_2), .IN1(1'b0), .IN2(~na318_2), .IN3(na233_1), .IN4(na218_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x42y120     80'h00_0018_00_0000_0C88_83FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_1 ( .OUT(na39_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na345_2), .IN7(na344_2), .IN8(na36_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x40y118     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a40_4 ( .OUT(na40_2), .IN1(~na258_2), .IN2(1'b0), .IN3(~na317_2), .IN4(na218_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x34y123     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a42_1 ( .OUT(na42_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(na148_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x36y119     80'h00_0018_00_0000_0888_EF53
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a43_1 ( .OUT(na43_1), .IN1(1'b0), .IN2(~na318_2), .IN3(~na44_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na234_1), .IN8(na218_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x38y121     80'h00_0078_00_0000_0C88_C841
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a44_1 ( .OUT(na44_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na214_2), .IN6(na345_2), .IN7(1'b1), .IN8(na218_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a44_4 ( .OUT(na44_2), .IN1(~na214_2), .IN2(~na148_1), .IN3(~na346_2), .IN4(na218_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x35y121     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a45_4 ( .OUT(na45_2), .IN1(na214_2), .IN2(~na148_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x39y118     80'h00_0060_00_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a46_4 ( .OUT(na46_2), .IN1(~na262_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x38y123     80'h00_0018_00_0040_0ACC_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a47_1 ( .OUT(na47_1), .IN1(1'b1), .IN2(na148_1), .IN3(1'b1), .IN4(~na335_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na341_2), .IN8(~na218_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x35y119     80'h00_0018_00_0000_0C88_E3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a48_1 ( .OUT(na48_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na318_2), .IN7(na235_1), .IN8(na218_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x38y117     80'h00_0018_00_0000_0888_5FD5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a49_1 ( .OUT(na49_1), .IN1(~na321_2), .IN2(1'b0), .IN3(~na236_1), .IN4(na218_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na44_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x31y122     80'h00_0060_00_0000_0C08_FFE5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a51_4 ( .OUT(na51_2), .IN1(~na321_2), .IN2(1'b0), .IN3(na237_1), .IN4(na218_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y119     80'h00_0018_00_0040_0AA2_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a52_1 ( .OUT(na52_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na218_1), .IN5(1'b0), .IN6(~na266_2), .IN7(1'b0), .IN8(na238_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x36y120     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a53_4 ( .OUT(na53_2), .IN1(~na214_2), .IN2(na148_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x40y120     80'h00_0018_00_0000_0888_EF55
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a54_1 ( .OUT(na54_1), .IN1(~na55_1), .IN2(1'b0), .IN3(~na44_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na239_1), .IN8(na218_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y121     80'h00_0018_00_0000_0C88_83FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na345_2), .IN7(na344_2), .IN8(na53_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x32y123     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a56_4 ( .OUT(na56_2), .IN1(~na55_1), .IN2(1'b0), .IN3(~na240_1), .IN4(na218_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x33y117     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a57_1 ( .OUT(na57_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na322_2), .IN6(1'b0), .IN7(~na241_1), .IN8(na218_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x39y118     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a58_1 ( .OUT(na58_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na321_2), .IN6(1'b0), .IN7(~na242_1), .IN8(na218_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x42y119     80'h00_0018_00_0000_0888_5FD3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a59_1 ( .OUT(na59_1), .IN1(1'b0), .IN2(~na318_2), .IN3(~na243_1), .IN4(na218_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na44_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x39y114     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a60_4 ( .OUT(na60_2), .IN1(1'b1), .IN2(~na32_2), .IN3(na250_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x40y121     80'h00_EA00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a61_4 ( .OUT(na61_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na49_1), .IN4(na21_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a61_5 ( .OUT(na61_2), .CLK(na163_1), .EN(na80_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na61_2_i) );
// C_AND/D///      x41y112     80'h00_EA00_00_0000_0C88_24FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a62_1 ( .OUT(na62_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na78_2), .IN6(na24_1), .IN7(na308_2), .IN8(~na29_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a62_2 ( .OUT(na62_1), .CLK(na163_1), .EN(na75_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na62_1_i) );
// C_ORAND////      x43y119     80'h00_0018_00_0000_0888_DCBE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a63_1 ( .OUT(na63_1), .IN1(na65_1), .IN2(na67_1), .IN3(na328_2), .IN4(~na21_1), .IN5(1'b0), .IN6(na70_1), .IN7(~na22_1),
                    .IN8(na327_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x37y113     80'h00_0018_00_0040_0C79_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a65_1 ( .OUT(na65_1), .IN1(~na28_1), .IN2(1'b1), .IN3(1'b1), .IN4(na309_2), .IN5(1'b1), .IN6(na24_1), .IN7(1'b1), .IN8(na29_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x43y121     80'h00_0078_00_0000_0C88_CAC3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a66_1 ( .OUT(na66_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na78_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a66_4 ( .OUT(na66_2), .IN1(1'b1), .IN2(~na24_1), .IN3(1'b1), .IN4(na12_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x41y118     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_1 ( .OUT(na67_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na312_2), .IN6(~na32_1), .IN7(~na31_1), .IN8(~na33_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x35y114     80'h00_0018_00_0040_0A36_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a70_1 ( .OUT(na70_1), .IN1(na28_1), .IN2(1'b1), .IN3(1'b1), .IN4(na29_2), .IN5(na273_1), .IN6(~na24_1), .IN7(1'b1), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x30y115     80'h00_EA00_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a71_1 ( .OUT(na71_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na24_1), .IN7(na27_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a71_2 ( .OUT(na71_1), .CLK(na163_1), .EN(na91_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na71_1_i) );
// C_ORAND*/DST///      x42y121     80'h20_BE00_00_0000_0788_F5DD
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a72_1 ( .OUT(na72_1_i), .IN1(~na66_1), .IN2(na19_1), .IN3(~na72_1), .IN4(na2_2), .IN5(~na66_2), .IN6(1'b0), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'bX_0100_0000)) 
           _a72_2 ( .OUT(na72_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na72_1_i) );
// C_///AND/D      x40y115     80'h00_EE00_80_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a74_4 ( .OUT(na74_2_i), .IN1(~na66_2), .IN2(na275_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a74_5 ( .OUT(na74_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na74_2_i) );
// C_MX4b////      x35y122     80'h00_0018_00_0040_0A51_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1), .IN1(1'b1), .IN2(na311_2), .IN3(na307_2), .IN4(1'b1), .IN5(~na28_1), .IN6(1'b0), .IN7(na276_1), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x30y118     80'h00_EE00_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a77_1 ( .OUT(na77_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na66_2), .IN6(1'b1), .IN7(na278_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a77_2 ( .OUT(na77_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na77_1_i) );
// C_///ORAND/D      x41y119     80'h00_EE00_80_0000_0C08_FFE5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a78_4 ( .OUT(na78_2_i), .IN1(~na66_2), .IN2(1'b0), .IN3(na79_2), .IN4(na280_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a78_5 ( .OUT(na78_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_2_i) );
// C_///ORAND/      x36y117     80'h00_0060_00_0000_0C08_FFBA
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a79_4 ( .OUT(na79_2), .IN1(na78_2), .IN2(1'b0), .IN3(na27_1), .IN4(~na2_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x31y121     80'h00_0018_00_0000_0888_ABBE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1), .IN1(na65_1), .IN2(na67_1), .IN3(na328_2), .IN4(~na21_1), .IN5(na66_1), .IN6(~na306_2), .IN7(na22_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x37y114     80'h00_0018_00_0000_0888_FCE3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a81_1 ( .OUT(na81_1), .IN1(1'b0), .IN2(~na333_2), .IN3(na74_2), .IN4(na83_1), .IN5(1'b0), .IN6(na85_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x40y112     80'h00_0018_00_0040_0AB7_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a83_1 ( .OUT(na83_1), .IN1(~na28_1), .IN2(1'b1), .IN3(1'b1), .IN4(na29_2), .IN5(~na282_1), .IN6(~na24_1), .IN7(1'b1), .IN8(na332_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x38y112     80'h00_0060_00_0000_0C08_FFA2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a84_4 ( .OUT(na84_2), .IN1(na66_1), .IN2(~na67_1), .IN3(na22_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x33y112     80'h00_0018_00_0040_0A68_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a85_1 ( .OUT(na85_1), .IN1(~na28_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2_2), .IN5(1'b0), .IN6(na283_1), .IN7(na347_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x31y115     80'h00_0018_00_0040_0A9D_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a88_1 ( .OUT(na88_1), .IN1(1'b1), .IN2(~na301_2), .IN3(1'b1), .IN4(~na309_2), .IN5(~na286_1), .IN6(1'b0), .IN7(1'b1), .IN8(~na29_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x31y123     80'h00_0018_00_0000_0C88_2CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na301_2), .IN7(na71_1), .IN8(~na272_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x32y114     80'h00_0018_00_0040_0AC8_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1), .IN1(na66_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na84_2), .IN5(1'b0), .IN6(1'b0), .IN7(na326_2), .IN8(~na272_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x31y120     80'h00_0018_00_0040_0AC8_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a91_1 ( .OUT(na91_1), .IN1(na66_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na92_2), .IN8(~na272_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x32y117     80'h00_0060_00_0000_0C08_FF82
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a92_4 ( .OUT(na92_2), .IN1(na329_2), .IN2(~na24_1), .IN3(na27_1), .IN4(na2_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x37y117     80'h00_0060_00_0000_0C08_FFE3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a93_4 ( .OUT(na93_2), .IN1(1'b0), .IN2(~na94_1), .IN3(na72_1), .IN4(na13_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x39y124     80'h00_0018_00_0040_0A9A_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a94_1 ( .OUT(na94_1), .IN1(1'b1), .IN2(~na301_2), .IN3(~na307_2), .IN4(1'b1), .IN5(na288_2), .IN6(1'b1), .IN7(1'b0), .IN8(~na12_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x37y124     80'h00_0018_00_0040_0A9B_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a102_1 ( .OUT(na102_1), .IN1(na150_1), .IN2(1'b1), .IN3(1'b1), .IN4(na218_2), .IN5(~na289_1), .IN6(1'b1), .IN7(1'b0), .IN8(~na218_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x36y124     80'h00_0018_00_0040_0A9A_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_1 ( .OUT(na103_1), .IN1(1'b1), .IN2(~na148_1), .IN3(1'b1), .IN4(na218_1), .IN5(na290_2), .IN6(1'b1), .IN7(1'b0), .IN8(~na218_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x35y118     80'h00_0018_00_0000_0C66_CBFF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a104_1 ( .OUT(na104_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na214_2), .IN6(na102_1), .IN7(1'b1), .IN8(~na103_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x32y116     80'h00_0018_00_0040_0C61_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a105_1 ( .OUT(na105_1), .IN1(na292_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b0), .IN5(na150_1), .IN6(1'b1), .IN7(1'b1), .IN8(na36_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x38y124     80'h00_0018_00_0040_0AA2_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a106_1 ( .OUT(na106_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na218_1), .IN5(1'b0), .IN6(~na37_2), .IN7(1'b0), .IN8(na105_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x40y117     80'h00_0018_00_0040_0C94_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a107_1 ( .OUT(na107_1), .IN1(1'b1), .IN2(1'b0), .IN3(na294_2), .IN4(1'b1), .IN5(na28_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na29_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x42y118     80'h00_0018_00_0000_0888_3A15
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a108_1 ( .OUT(na108_1), .IN1(~na295_2), .IN2(1'b1), .IN3(~na26_1), .IN4(~na284_2), .IN5(na88_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na284_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x32y119     80'h00_0078_00_0020_0C66_CCCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a110_1 ( .OUT(na110_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na148_1), .IN7(1'b1), .IN8(na342_2),
                     .CINX(1'b0), .CINY1(na116_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a110_4 ( .OUT(na110_2), .COUTY1(na110_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na218_2), .IN5(1'b1), .IN6(na148_1), .IN7(1'b1),
                     .IN8(na342_2), .CINX(1'b0), .CINY1(na116_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x32y120     80'h00_0078_00_0020_0C66_FACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a112_1 ( .OUT(na112_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na150_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na110_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a112_4 ( .OUT(na112_2), .COUTY1(na112_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na218_1), .IN5(na150_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na110_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x32y121     80'h00_0078_00_0020_0C66_FCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a114_1 ( .OUT(na114_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na152_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na112_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a114_4 ( .OUT(na114_2), .COUTY1(na114_4), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(na220_1), .IN5(1'b1), .IN6(na152_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na112_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x32y118     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a116_2 ( .OUT(na116_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a116_6 ( .COUTY1(na116_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na116_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x29y119     80'h00_0078_00_0020_0C66_CAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a117_1 ( .OUT(na117_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na8_2), .IN6(1'b1), .IN7(1'b1), .IN8(na302_2),
                     .CINX(1'b0), .CINY1(na123_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a117_4 ( .OUT(na117_2), .COUTY1(na117_4), .IN1(1'b0), .IN2(1'b0), .IN3(na5_1), .IN4(1'b1), .IN5(na8_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na302_2), .CINX(1'b0), .CINY1(na123_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x29y120     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a119_1 ( .OUT(na119_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na5_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na117_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a119_4 ( .OUT(na119_2), .COUTY1(na119_4), .IN1(1'b1), .IN2(na4_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na5_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na117_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x29y121     80'h00_0078_00_0020_0C66_0AC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a121_1 ( .OUT(na121_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na8_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na119_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a121_4 ( .OUT(na121_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na9_2), .IN5(na8_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na119_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x29y118     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a123_2 ( .OUT(na123_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a123_6 ( .COUTY1(na123_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na123_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x34y115     80'h00_EE60_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a125_1 ( .OUT(na125_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na125_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na146_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a125_2 ( .OUT(na125_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na125_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a125_4 ( .OUT(na125_2), .COUTY1(na125_4), .IN1(1'b0), .IN2(1'b0), .IN3(na175_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na125_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na146_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y116     80'h00_EE60_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a127_1 ( .OUT(na127_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na127_1),
                     .CINX(1'b0), .CINY1(na125_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a127_2 ( .OUT(na127_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na127_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a127_4 ( .OUT(na127_2), .COUTY1(na127_4), .IN1(na177_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na127_1), .CINX(1'b0), .CINY1(na125_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y117     80'h00_EE60_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a129_1 ( .OUT(na129_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na129_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na127_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a129_2 ( .OUT(na129_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na129_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a129_4 ( .OUT(na129_2), .COUTY1(na129_4), .IN1(1'b1), .IN2(na179_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na129_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na127_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y118     80'h00_EE60_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a131_1 ( .OUT(na131_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na131_1),
                     .CINX(1'b0), .CINY1(na129_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a131_2 ( .OUT(na131_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na131_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a131_4 ( .OUT(na131_2), .COUTY1(na131_4), .IN1(1'b0), .IN2(1'b0), .IN3(na181_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na131_1), .CINX(1'b0), .CINY1(na129_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y119     80'h00_EE60_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a133_1 ( .OUT(na133_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na133_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na131_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a133_2 ( .OUT(na133_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na133_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a133_4 ( .OUT(na133_2), .COUTY1(na133_4), .IN1(na183_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na133_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na131_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y110     80'h00_EE60_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a134_1 ( .OUT(na134_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na165_2), .IN6(1'b1), .IN7(1'b1), .IN8(na134_1),
                     .CINX(1'b0), .CINY1(na147_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a134_2 ( .OUT(na134_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na134_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a134_4 ( .OUT(na134_2), .COUTY1(na134_4), .IN1(na165_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na165_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na134_1), .CINX(1'b0), .CINY1(na147_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y120     80'h00_EE60_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a136_1 ( .OUT(na136_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na136_1),
                     .CINX(1'b0), .CINY1(na133_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a136_2 ( .OUT(na136_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na136_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a136_4 ( .OUT(na136_2), .COUTY1(na136_4), .IN1(1'b0), .IN2(1'b0), .IN3(na185_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na136_1), .CINX(1'b0), .CINY1(na133_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF/D///      x34y121     80'h00_EE00_00_0010_0666_00A0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a138_1 ( .OUT(na138_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na138_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na136_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a138_2 ( .OUT(na138_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na138_1_i) );
// C_ADDF2/D//ADDF2/      x34y111     80'h00_EE60_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a140_1 ( .OUT(na140_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na140_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na134_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a140_2 ( .OUT(na140_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na140_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a140_4 ( .OUT(na140_2), .COUTY1(na140_4), .IN1(1'b0), .IN2(1'b0), .IN3(na167_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na140_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na134_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y112     80'h00_EE60_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a142_1 ( .OUT(na142_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na142_1),
                     .CINX(1'b0), .CINY1(na140_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a142_2 ( .OUT(na142_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na142_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a142_4 ( .OUT(na142_2), .COUTY1(na142_4), .IN1(1'b0), .IN2(1'b0), .IN3(na169_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na142_1), .CINX(1'b0), .CINY1(na140_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y113     80'h00_EE60_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a144_1 ( .OUT(na144_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na144_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na142_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a144_2 ( .OUT(na144_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na144_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a144_4 ( .OUT(na144_2), .COUTY1(na144_4), .IN1(1'b0), .IN2(1'b0), .IN3(na171_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na144_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na142_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x34y114     80'h00_EE60_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a146_1 ( .OUT(na146_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na146_1),
                     .CINX(1'b0), .CINY1(na144_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a146_2 ( .OUT(na146_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na146_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a146_4 ( .OUT(na146_2), .COUTY1(na146_4), .IN1(na173_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na146_1), .CINX(1'b0), .CINY1(na144_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x34y109     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a147_2 ( .OUT(na147_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a147_6 ( .COUTY1(na147_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na147_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x33y122     80'h00_EA60_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a148_1 ( .OUT(na148_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na148_1), .IN7(1'b1), .IN8(na342_2),
                     .CINX(1'b0), .CINY1(na154_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a148_2 ( .OUT(na148_1), .CLK(na163_1), .EN(na89_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na148_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a148_4 ( .OUT(na148_2), .COUTY1(na148_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na218_2), .IN5(1'b1), .IN6(na148_1), .IN7(1'b1),
                     .IN8(na342_2), .CINX(1'b0), .CINY1(na154_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x33y123     80'h00_EA60_00_0020_0C66_0AC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a150_1 ( .OUT(na150_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na150_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na148_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a150_2 ( .OUT(na150_1), .CLK(na163_1), .EN(na89_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na150_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a150_4 ( .OUT(na150_2), .COUTY1(na150_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na218_1), .IN5(na150_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na148_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x33y124     80'h00_EA60_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a152_1 ( .OUT(na152_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na152_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na150_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a152_2 ( .OUT(na152_1), .CLK(na163_1), .EN(na89_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na152_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a152_4 ( .OUT(na152_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na220_1), .IN5(1'b1), .IN6(na152_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na150_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x33y121     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a154_2 ( .OUT(na154_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a154_6 ( .COUTY1(na154_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na154_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x41y115     80'h00_0078_00_0020_0C66_ACFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a155_1 ( .OUT(na155_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na32_2), .IN7(na31_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na158_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a155_4 ( .OUT(na155_2), .COUTY1(na155_4), .IN1(1'b1), .IN2(na32_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na32_2), .IN7(na31_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na158_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x41y116     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a157_1 ( .OUT(na157_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na33_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na155_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x41y114     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a158_2 ( .OUT(na158_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a158_6 ( .COUTY1(na158_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na158_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x38y114     80'h00_0078_00_0020_0C66_ACFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a159_1 ( .OUT(na159_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na32_2), .IN7(na31_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na260_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a159_4 ( .OUT(na159_2), .COUTY1(na159_4), .IN1(1'b1), .IN2(na32_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na32_2), .IN7(na31_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na260_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x38y115     80'h00_0018_00_0010_0666_00CF
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a161_1 ( .OUT(na161_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na33_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na159_4), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0000_0010)) 
           _a163 ( .GLB0(na163_1), .GLB1(_d3), .GLB2(_d4), .GLB3(_d5), .CLK_FB0(_d6), .CLK_FB1(_d7), .CLK_FB2(_d8), .CLK_FB3(_d9),
                   .CLK0_0(1'b0), .CLK0_90(1'b0), .CLK0_180(1'b0), .CLK0_270(1'b0), .CLK0_BYP(na1_1), .CLK1_0(1'b0), .CLK1_90(1'b0),
                   .CLK1_180(1'b0), .CLK1_270(1'b0), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0), .CLK2_270(1'b0),
                   .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0), .USR_GLB0(1'b0),
                   .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0), .USR_FB3(1'b0) );
// C_AND/D//AND/D      x29y109     80'h00_EE00_80_0000_0C88_CFF5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a165_1 ( .OUT(na165_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na134_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a165_2 ( .OUT(na165_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na165_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a165_4 ( .OUT(na165_2_i), .IN1(~na165_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a165_5 ( .OUT(na165_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na165_2_i) );
// C_///AND/D      x32y109     80'h00_EE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a167_4 ( .OUT(na167_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na140_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a167_5 ( .OUT(na167_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na167_2_i) );
// C_AND/D///      x32y109     80'h00_EE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a169_1 ( .OUT(na169_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na142_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a169_2 ( .OUT(na169_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na169_1_i) );
// C_///AND/D      x32y111     80'h00_EE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a171_4 ( .OUT(na171_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na144_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a171_5 ( .OUT(na171_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na171_2_i) );
// C_AND/D///      x33y113     80'h00_EE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a173_1 ( .OUT(na173_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na146_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a173_2 ( .OUT(na173_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na173_1_i) );
// C_///AND/D      x30y113     80'h00_EE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a175_4 ( .OUT(na175_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na125_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a175_5 ( .OUT(na175_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na175_2_i) );
// C_///AND/D      x33y115     80'h00_EE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a177_4 ( .OUT(na177_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na127_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a177_5 ( .OUT(na177_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na177_2_i) );
// C_AND/D///      x33y118     80'h00_EE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a179_1 ( .OUT(na179_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na129_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a179_2 ( .OUT(na179_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na179_1_i) );
// C_///AND/D      x30y117     80'h00_EE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a181_4 ( .OUT(na181_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na131_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a181_5 ( .OUT(na181_2), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na181_2_i) );
// C_AND/D///      x35y117     80'h00_EE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a183_1 ( .OUT(na183_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na133_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a183_2 ( .OUT(na183_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na183_1_i) );
// C_AND/D///      x30y119     80'h00_EE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a185_1 ( .OUT(na185_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na136_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a185_2 ( .OUT(na185_1), .CLK(na163_1), .EN(1'b1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na185_1_i) );
// C_///AND/D      x31y123     80'h00_EA00_80_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a214_4 ( .OUT(na214_2_i), .IN1(~na214_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a214_5 ( .OUT(na214_2), .CLK(na163_1), .EN(na89_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na214_2_i) );
// C_AND/D//AND/D      x38y120     80'h00_EA00_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a218_1 ( .OUT(na218_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na150_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a218_2 ( .OUT(na218_1), .CLK(na163_1), .EN(na89_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na218_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a218_4 ( .OUT(na218_2_i), .IN1(1'b1), .IN2(na148_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a218_5 ( .OUT(na218_2), .CLK(na163_1), .EN(na89_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na218_2_i) );
// C_AND/D///      x30y124     80'h00_EA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a220_1 ( .OUT(na220_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na152_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a220_2 ( .OUT(na220_1), .CLK(na163_1), .EN(na89_1), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na220_1_i) );
// C_MX4b////      x35y112     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a222_1 ( .OUT(na222_1), .IN1(1'b1), .IN2(na32_2), .IN3(1'b1), .IN4(na159_1), .IN5(na38_2), .IN6(na104_1), .IN7(na43_1), .IN8(na40_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x35y115     80'h00_0018_00_0040_0AF4_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a223_1 ( .OUT(na223_1), .IN1(1'b1), .IN2(na32_2), .IN3(1'b1), .IN4(na159_1), .IN5(na48_1), .IN6(na46_2), .IN7(~na49_1), .IN8(na106_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x42y116     80'h00_0018_00_0040_0AF4_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a224_1 ( .OUT(na224_1), .IN1(1'b1), .IN2(na32_2), .IN3(1'b1), .IN4(na159_1), .IN5(na52_1), .IN6(na51_2), .IN7(~na56_2), .IN8(na54_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x32y115     80'h00_0018_00_0040_0A77_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a225_1 ( .OUT(na225_1), .IN1(1'b1), .IN2(~na32_2), .IN3(1'b1), .IN4(na159_1), .IN5(~na57_1), .IN6(~na58_1), .IN7(~na59_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x37y115     80'h00_0018_00_0040_0AF0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a226_1 ( .OUT(na226_1), .IN1(1'b1), .IN2(~na339_2), .IN3(na161_1), .IN4(1'b1), .IN5(na223_1), .IN6(na222_1), .IN7(na225_1),
                     .IN8(na224_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x39y121     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a227_1 ( .OUT(na227_1), .IN1(1'b1), .IN2(na32_2), .IN3(1'b1), .IN4(na336_2), .IN5(na38_2), .IN6(na104_1), .IN7(na43_1), .IN8(na40_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x39y116     80'h00_0018_00_0040_0AF4_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a228_1 ( .OUT(na228_1), .IN1(1'b1), .IN2(na32_2), .IN3(1'b1), .IN4(na336_2), .IN5(na48_1), .IN6(na46_2), .IN7(~na49_1), .IN8(na106_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x40y123     80'h00_0018_00_0040_0AF4_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a229_1 ( .OUT(na229_1), .IN1(1'b1), .IN2(na32_2), .IN3(1'b1), .IN4(na336_2), .IN5(na52_1), .IN6(na51_2), .IN7(~na56_2), .IN8(na54_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x38y122     80'h00_0018_00_0040_0A77_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a230_1 ( .OUT(na230_1), .IN1(1'b1), .IN2(~na32_2), .IN3(1'b1), .IN4(na336_2), .IN5(~na57_1), .IN6(~na58_1), .IN7(~na59_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x44y121     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a231_1 ( .OUT(na231_1), .IN1(na155_2), .IN2(1'b1), .IN3(1'b1), .IN4(na337_2), .IN5(na227_1), .IN6(na228_1), .IN7(na229_1),
                     .IN8(na230_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x43y114     80'h00_0018_00_0040_0AE0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a232_1 ( .OUT(na232_1), .IN1(1'b1), .IN2(na338_2), .IN3(1'b1), .IN4(na159_2), .IN5(1'b0), .IN6(na60_2), .IN7(na325_2), .IN8(na14_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x36y123     80'h00_0018_00_0040_0AF1_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a233_1 ( .OUT(na233_1), .IN1(~na150_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na218_2), .IN5(~na315_2), .IN6(na324_2), .IN7(na42_1),
                     .IN8(na35_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x36y121     80'h00_0018_00_0040_0AD2_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a234_1 ( .OUT(na234_1), .IN1(~na150_1), .IN2(1'b1), .IN3(1'b1), .IN4(na218_2), .IN5(na45_2), .IN6(1'b1), .IN7(na42_1), .IN8(na36_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x28y119     80'h00_0018_00_0040_0AD2_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a235_1 ( .OUT(na235_1), .IN1(1'b1), .IN2(~na345_2), .IN3(1'b1), .IN4(na335_2), .IN5(na313_2), .IN6(1'b1), .IN7(na42_1), .IN8(na35_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x38y119     80'h00_0018_00_0040_0AEB_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a236_1 ( .OUT(na236_1), .IN1(~na150_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na218_2), .IN5(1'b1), .IN6(~na148_1), .IN7(na42_1),
                     .IN8(~na320_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x36y125     80'h00_0018_00_0040_0AFD_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a237_1 ( .OUT(na237_1), .IN1(na150_1), .IN2(1'b1), .IN3(1'b1), .IN4(na218_2), .IN5(~na214_2), .IN6(na340_2), .IN7(~na42_1),
                     .IN8(~na36_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x34y124     80'h00_0018_00_0040_0AF8_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a238_1 ( .OUT(na238_1), .IN1(1'b1), .IN2(~na345_2), .IN3(1'b1), .IN4(~na335_2), .IN5(na45_2), .IN6(na148_1), .IN7(na334_2),
                     .IN8(~na53_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x34y125     80'h00_0018_00_0040_0AD9_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a239_1 ( .OUT(na239_1), .IN1(1'b1), .IN2(~na345_2), .IN3(1'b1), .IN4(~na335_2), .IN5(~na45_2), .IN6(1'b0), .IN7(na42_1),
                     .IN8(~na323_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x34y127     80'h00_0018_00_0040_0AF7_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a240_1 ( .OUT(na240_1), .IN1(~na150_1), .IN2(1'b1), .IN3(1'b1), .IN4(na218_2), .IN5(~na45_2), .IN6(~na316_2), .IN7(~na42_1),
                     .IN8(na35_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x38y125     80'h00_0018_00_0040_0A36_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a241_1 ( .OUT(na241_1), .IN1(na150_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na218_2), .IN5(na214_2), .IN6(~na314_2), .IN7(1'b1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x36y127     80'h00_0018_00_0040_0AF0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a242_1 ( .OUT(na242_1), .IN1(~na150_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na218_2), .IN5(na313_2), .IN6(na148_1), .IN7(na42_1),
                     .IN8(na36_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x40y125     80'h00_0018_00_0040_0AB2_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a243_1 ( .OUT(na243_1), .IN1(na150_1), .IN2(1'b1), .IN3(1'b1), .IN4(na218_2), .IN5(na319_2), .IN6(~na148_1), .IN7(1'b0),
                     .IN8(na36_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a244 ( .Y(na244_1), .I(areset_n) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a245 ( .Y(na245_1), .I(clk_10MHz) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a246 ( .O(led), .A(na296_10) );
CPE_IOBF   #(.BUF_CFG (72'h00000100010006091C)) 
           _a247 ( .Y(_d10), .O(i2c_scl), .A(na297_10), .EN(na298_10) );
CPE_IOBF   #(.BUF_CFG (72'h00000100010006091C)) 
           _a248 ( .Y(na248_1), .O(i2c_sda), .A(na299_10), .EN(na300_10) );
// C_AND///AND/      x43y120     80'h00_0078_00_0000_0C88_F4CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a249_1 ( .OUT(na249_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na65_1), .IN6(na232_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a249_4 ( .OUT(na249_2), .IN1(1'b1), .IN2(na24_1), .IN3(1'b1), .IN4(na29_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x38y111     80'h00_EA00_80_0000_0C08_FFFF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a250_4 ( .OUT(na250_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a250_5 ( .OUT(na250_2), .CLK(na163_1), .EN(na66_2), .SR(na244_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na250_2_i) );
// C_///AND/      x40y114     80'h00_0060_00_0000_0C08_FF15
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a252_4 ( .OUT(na252_2), .IN1(~na305_2), .IN2(1'b1), .IN3(~na26_1), .IN4(~na21_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y120     80'h00_0018_00_0000_0C88_51FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a253_1 ( .OUT(na253_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na305_2), .IN6(~na23_2), .IN7(~na26_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y112     80'h00_0018_00_0000_0C88_2CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a254_1 ( .OUT(na254_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na24_1), .IN7(na22_2), .IN8(~na29_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x36y118     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a256_1 ( .OUT(na256_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na78_2), .IN6(1'b1), .IN7(~na161_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y123     80'h00_0060_00_0000_0C08_FFC2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a258_4 ( .OUT(na258_2), .IN1(na150_1), .IN2(~na343_2), .IN3(1'b1), .IN4(na259_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x34y122     80'h00_0060_00_0000_0C0E_FF75
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a259_4 ( .OUT(na259_2), .IN1(~na150_1), .IN2(1'b0), .IN3(~na42_1), .IN4(~na218_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x38y113     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a260_2 ( .OUT(na260_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a260_6 ( .COUTY1(na260_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na260_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x33y117     80'h00_0060_00_0000_0C08_FF43
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a262_4 ( .OUT(na262_2), .IN1(1'b1), .IN2(~na343_2), .IN3(~na47_1), .IN4(na259_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x35y120     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a266_4 ( .OUT(na266_2), .IN1(na214_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na218_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x32y122     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a272_1 ( .OUT(na272_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0), .CINX(1'b0),
                     .CINY1(na114_4), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y115     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a273_1 ( .OUT(na273_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na24_1), .IN7(1'b1), .IN8(~na272_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x41y122     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a275_1 ( .OUT(na275_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na2_2), .IN5(na331_2), .IN6(1'b0), .IN7(na74_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x42y113     80'h00_0018_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a276_1 ( .OUT(na276_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na28_1), .IN6(1'b1), .IN7(na277_1), .IN8(na2_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y111     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a277_1 ( .OUT(na277_1), .IN1(1'b1), .IN2(na330_2), .IN3(1'b0), .IN4(1'b0), .IN5(na78_2), .IN6(~na248_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x28y113     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a278_1 ( .OUT(na278_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na2_2), .IN5(na331_2), .IN6(1'b0), .IN7(na72_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x36y112     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a280_1 ( .OUT(na280_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na74_2), .IN8(na2_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x41y121     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a282_1 ( .OUT(na282_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na78_2), .IN6(~na24_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x31y114     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a283_1 ( .OUT(na283_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na24_1), .IN7(1'b1), .IN8(~na29_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x36y114     80'h00_0078_00_0000_0C88_AC3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_1 ( .OUT(na284_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na67_1), .IN7(na22_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a284_4 ( .OUT(na284_2), .IN1(1'b1), .IN2(na24_1), .IN3(1'b1), .IN4(~na2_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x39y117     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a286_1 ( .OUT(na286_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na74_2), .IN8(na29_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x41y113     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a288_4 ( .OUT(na288_2), .IN1(~na78_2), .IN2(1'b1), .IN3(1'b1), .IN4(na12_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x31y125     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a289_1 ( .OUT(na289_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na148_1), .IN7(1'b1), .IN8(~na218_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x35y123     80'h00_0060_00_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a290_4 ( .OUT(na290_2), .IN1(~na150_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na218_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x31y119     80'h00_0060_00_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a292_4 ( .OUT(na292_2), .IN1(~na214_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na218_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x42y113     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a294_4 ( .OUT(na294_2), .IN1(1'b1), .IN2(na24_1), .IN3(1'b1), .IN4(~na77_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x35y111     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a295_4 ( .OUT(na295_2), .IN1(~na78_2), .IN2(1'b1), .IN3(na107_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x1y95     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a296_4 ( .OUT(na296_2), .IN1(1'b1), .IN2(1'b1), .IN3(na138_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a296_6 ( .RAM_O2(na296_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na296_2), .COMP_OUT(1'b0) );
// C_///AND/      x57y128     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a297_4 ( .OUT(na297_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a297_6 ( .RAM_O2(na297_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na297_2), .COMP_OUT(1'b0) );
// C_///AND/      x58y128     80'h08_0060_00_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a298_4 ( .OUT(na298_2), .IN1(1'b1), .IN2(~na10_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a298_6 ( .RAM_O2(na298_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na298_2), .COMP_OUT(1'b0) );
// C_///AND/      x59y128     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a299_4 ( .OUT(na299_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a299_6 ( .RAM_O2(na299_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na299_2), .COMP_OUT(1'b0) );
// C_///AND/      x60y128     80'h08_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a300_4 ( .OUT(na300_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na15_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a300_6 ( .RAM_O2(na300_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na300_2), .COMP_OUT(1'b0) );
// C_////Bridge      x33y118     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a301_5 ( .OUT(na301_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y118     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a302_5 ( .OUT(na302_2), .IN1(1'b0), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y115     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a303_5 ( .OUT(na303_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na12_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y115     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a304_5 ( .OUT(na304_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na19_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y117     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a305_5 ( .OUT(na305_2), .IN1(1'b0), .IN2(1'b0), .IN3(na22_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y120     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a306_5 ( .OUT(na306_2), .IN1(1'b0), .IN2(1'b0), .IN3(na22_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y119     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a307_5 ( .OUT(na307_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na24_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y111     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a308_5 ( .OUT(na308_2), .IN1(na28_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y112     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a309_5 ( .OUT(na309_2), .IN1(na28_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a310_5 ( .OUT(na310_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na29_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y120     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a311_5 ( .OUT(na311_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na29_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y115     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a312_5 ( .OUT(na312_2), .IN1(1'b0), .IN2(na32_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y121     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a313_5 ( .OUT(na313_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na35_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y126     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a314_5 ( .OUT(na314_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na35_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y123     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a315_5 ( .OUT(na315_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na36_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y128     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a316_5 ( .OUT(na316_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na36_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a317_5 ( .OUT(na317_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na36_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y120     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a318_5 ( .OUT(na318_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na39_1) );
// C_////Bridge      x41y125     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a319_5 ( .OUT(na319_2), .IN1(1'b0), .IN2(1'b0), .IN3(na42_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y122     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a320_5 ( .OUT(na320_2), .IN1(1'b0), .IN2(1'b0), .IN3(na42_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y119     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a321_5 ( .OUT(na321_2), .IN1(1'b0), .IN2(1'b0), .IN3(na44_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y115     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a322_5 ( .OUT(na322_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na44_2), .IN8(1'b0) );
// C_////Bridge      x36y126     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a323_5 ( .OUT(na323_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na45_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y122     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a324_5 ( .OUT(na324_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na53_2) );
// C_////Bridge      x46y113     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a325_5 ( .OUT(na325_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na60_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x30y111     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a326_5 ( .OUT(na326_2), .IN1(na66_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y120     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a327_5 ( .OUT(na327_2), .IN1(na66_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y117     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a328_5 ( .OUT(na328_2), .IN1(1'b0), .IN2(na67_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y115     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a329_5 ( .OUT(na329_2), .IN1(1'b0), .IN2(1'b0), .IN3(na74_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y114     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a330_5 ( .OUT(na330_2), .IN1(1'b0), .IN2(1'b0), .IN3(na74_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y117     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a331_5 ( .OUT(na331_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na77_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y112     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a332_5 ( .OUT(na332_2), .IN1(na78_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y112     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a333_5 ( .OUT(na333_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na84_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y123     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a334_5 ( .OUT(na334_2), .IN1(1'b0), .IN2(na148_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y122     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a335_5 ( .OUT(na335_2), .IN1(na150_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y120     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a336_5 ( .OUT(na336_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na155_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y122     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a337_5 ( .OUT(na337_2), .IN1(1'b0), .IN2(na157_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y114     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a338_5 ( .OUT(na338_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na159_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y116     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a339_5 ( .OUT(na339_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na159_2) );
// C_////Bridge      x37y126     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a340_5 ( .OUT(na340_2), .IN1(na214_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y123     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a341_5 ( .OUT(na341_2), .IN1(na214_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x30y118     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a342_5 ( .OUT(na342_2), .IN1(na214_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y118     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a343_5 ( .OUT(na343_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na218_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y115     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a344_5 ( .OUT(na344_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na218_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y120     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a345_5 ( .OUT(na345_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na218_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y119     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a346_5 ( .OUT(na346_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na218_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y111     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a347_5 ( .OUT(na347_2), .IN1(1'b0), .IN2(na283_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
endmodule
