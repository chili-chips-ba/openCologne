//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 January 2025)
//  Compile Time: 2025-02-04 05:47:38
//  Program Run:  2025-03-16 11:26:34
//  Program Call: /home/tibrahimovic/0.git-repo/cc-toolchain-linux/bin/p_r/p_r -i net/FemtoRV32_synth.v -o FemtoRV32 -ccf /home/tibrahimovic/projects/femtorv32-quark-bicycle/3.build/../1.hw/constraints/constraints.ccf -cCP --verbose 
//  File Type:    Verilog

// Gatecount:   1516
module FemtoRV32 (clk , mem_rbusy , mem_rdata , mem_wbusy , reset ,
       mem_addr , mem_rstrb , mem_wdata , mem_wmask 
       ) ;

input  clk;
input  mem_rbusy;
input  [31:0]mem_rdata;
input  mem_wbusy;
input  reset;

output [31:0]mem_addr;
output mem_rstrb;
output [31:0]mem_wdata;
output [3:0]mem_wmask;



wire [31:0]mem_rdata;
wire [31:0]mem_addr;
wire [31:0]mem_wdata;
wire [3:0]mem_wmask;
wire clk;
wire na1_2;
wire na2_1;
wire na3_2;
wire na4_1;
wire na5_1;
wire na5_2;
wire na6_1;
wire na7_1;
wire na8_1;
wire na9_2;
wire reset;
wire na10_1;
wire na11_1;
wire na12_1;
wire na13_1;
wire na14_1;
wire na15_1;
wire na16_1;
wire na17_1;
wire na18_1;
wire na19_1;
wire na20_1;
wire na21_1;
wire na22_1;
wire na23_1;
wire na24_1;
wire na25_1;
wire na26_1;
wire na27_1;
wire na28_1;
wire na29_1;
wire na30_1;
wire na31_1;
wire na32_1;
wire na33_1;
wire na34_1;
wire na35_1;
wire na36_1;
wire na37_1;
wire na38_1;
wire na39_1;
wire na40_1;
wire na42_1;
wire na42_1_i;
wire na44_1;
wire na44_2;
wire na45_1;
wire na46_1;
wire na47_2;
wire na47_2_i;
wire na49_1;
wire na49_2;
wire na50_1;
wire na50_1_i;
wire na75_1;
wire na76_1;
wire na77_1;
wire na78_1;
wire na79_1;
wire na80_1;
wire na81_1;
wire na83_2;
wire na84_1;
wire na84_2;
wire na85_1;
wire na86_1;
wire na89_1;
wire na90_1;
wire na92_1;
wire na92_2;
wire na97_1;
wire na97_2;
wire na99_1;
wire na99_2;
wire na100_1;
wire na100_2;
wire na101_1;
wire na101_2;
wire na102_1;
wire na102_2;
wire na106_1;
wire na107_1;
wire na108_1;
wire na111_2;
wire na112_1;
wire na113_1;
wire na116_1;
wire na117_1;
wire na118_1;
wire na121_2;
wire na122_1;
wire na123_1;
wire na126_1;
wire na127_1;
wire na128_1;
wire na131_2;
wire na132_1;
wire na133_1;
wire na136_1;
wire na137_1;
wire na138_1;
wire na141_2;
wire na142_1;
wire na143_1;
wire na146_1;
wire na147_1;
wire na148_1;
wire na151_2;
wire na152_1;
wire na153_1;
wire na156_1;
wire na157_1;
wire na158_1;
wire na161_2;
wire na162_1;
wire na163_1;
wire na166_1;
wire na167_1;
wire na168_1;
wire na171_1;
wire na172_1;
wire na173_1;
wire na176_1;
wire na177_1;
wire na178_1;
wire na181_2;
wire na182_1;
wire na183_1;
wire na186_1;
wire na187_1;
wire na188_1;
wire na191_2;
wire na192_1;
wire na193_1;
wire na196_1;
wire na197_1;
wire na198_1;
wire na201_2;
wire na202_1;
wire na203_1;
wire na206_1;
wire na207_1;
wire na208_1;
wire na211_2;
wire na212_1;
wire na213_1;
wire na216_1;
wire na217_1;
wire na218_1;
wire na219_1;
wire na220_1;
wire na221_1;
wire na222_1;
wire na223_1;
wire na224_1;
wire na225_1;
wire na226_1;
wire na227_1;
wire na228_1;
wire na229_1;
wire na230_1;
wire na231_1;
wire na232_1;
wire na233_1;
wire na234_1;
wire na235_1;
wire na236_1;
wire na237_1;
wire na238_1;
wire na239_1;
wire na240_1;
wire na240_2;
wire na241_1;
wire na241_1_i;
wire na247_2;
wire na247_2_i;
wire na249_1;
wire na249_1_i;
wire na250_1;
wire na250_1_i;
wire na250_2;
wire na250_2_i;
wire na252_1;
wire na252_1_i;
wire na252_2;
wire na252_2_i;
wire na254_1;
wire na254_1_i;
wire na254_2;
wire na254_2_i;
wire na256_1;
wire na256_1_i;
wire na256_2;
wire na256_2_i;
wire na258_1;
wire na258_1_i;
wire na258_2;
wire na258_2_i;
wire na260_1;
wire na260_1_i;
wire na260_2;
wire na260_2_i;
wire na262_1;
wire na262_1_i;
wire na262_2;
wire na262_2_i;
wire na264_1;
wire na264_1_i;
wire na264_2;
wire na264_2_i;
wire na266_1;
wire na266_1_i;
wire na266_2;
wire na266_2_i;
wire na268_1;
wire na268_1_i;
wire na268_2;
wire na268_2_i;
wire na269_2;
wire na269_2_i;
wire na270_1;
wire na272_1;
wire na273_1;
wire na274_1;
wire na275_1;
wire na276_1;
wire na277_1;
wire na278_1;
wire na279_1;
wire na280_1;
wire na281_1;
wire na282_1;
wire na283_1;
wire na284_1;
wire na285_1;
wire na286_1;
wire na287_1;
wire na288_1;
wire na289_1;
wire na290_1;
wire na291_1;
wire na292_1;
wire na293_1;
wire na294_1;
wire na295_1;
wire na296_1;
wire na297_1;
wire na298_1;
wire na299_2;
wire na300_1;
wire na301_1;
wire na302_1;
wire na303_1;
wire na304_1;
wire na305_1;
wire na306_1;
wire na307_1;
wire na308_1;
wire na309_1;
wire na310_1;
wire na311_1;
wire na312_1;
wire na313_1;
wire na314_2;
wire na315_2;
wire na316_1;
wire na317_1;
wire na318_1;
wire na319_1;
wire na320_1;
wire na321_1;
wire na322_1;
wire na323_1;
wire na324_1;
wire na325_1;
wire na326_1;
wire na327_1;
wire na328_1;
wire na330_1;
wire na331_1;
wire na332_1;
wire na333_2;
wire na334_1;
wire na335_1;
wire na336_1;
wire na342_1;
wire na343_1;
wire na344_1;
wire na346_1;
wire na348_1;
wire na348_2;
wire na349_1;
wire na350_1;
wire na350_2;
wire na351_1;
wire na352_1;
wire na353_1;
wire na354_1;
wire na355_1;
wire na356_1;
wire na357_1;
wire na358_1;
wire na359_1;
wire na360_1;
wire na361_1;
wire na362_1;
wire na363_1;
wire na364_1;
wire na367_1;
wire na368_1;
wire na369_1;
wire na370_1;
wire na371_1;
wire na374_1;
wire na375_1;
wire na376_2;
wire na377_2;
wire na378_1;
wire na380_1;
wire na381_1;
wire na382_1;
wire na386_1;
wire na388_1;
wire na390_1;
wire na391_2;
wire na392_1;
wire na393_1;
wire na394_1;
wire na395_1;
wire na396_1;
wire na397_1;
wire na398_1;
wire na399_1;
wire na400_1;
wire na401_1;
wire na402_1;
wire na403_1;
wire na404_1;
wire na406_1;
wire na407_2;
wire na408_1;
wire na409_1;
wire na410_2;
wire na415_1;
wire na417_1;
wire na418_1;
wire na419_1;
wire na420_1;
wire na421_1;
wire na423_1;
wire na424_1;
wire na425_1;
wire na427_1;
wire na428_1;
wire na429_2;
wire na430_1;
wire na431_1;
wire na432_1;
wire na436_1;
wire na438_1;
wire na440_1;
wire na441_1;
wire na442_1;
wire na443_1;
wire na444_1;
wire na446_1;
wire na447_1;
wire na449_1;
wire na451_1;
wire na452_1;
wire na453_1;
wire na456_1;
wire na458_1;
wire na460_1;
wire na462_1;
wire na463_2;
wire na464_2;
wire na465_1;
wire na466_1;
wire na467_2;
wire na468_1;
wire na469_1;
wire na470_1;
wire na474_1;
wire na476_1;
wire na479_1;
wire na480_1;
wire na482_1;
wire na484_1;
wire na485_1;
wire na486_1;
wire na489_1;
wire na491_1;
wire na493_1;
wire na494_2;
wire na495_1;
wire na496_1;
wire na498_1;
wire na499_1;
wire na500_1;
wire na501_1;
wire na503_1;
wire na508_1;
wire na509_1;
wire na510_1;
wire na510_2;
wire na511_1;
wire na512_1;
wire na513_1;
wire na514_1;
wire na516_1;
wire na517_1;
wire na518_1;
wire na521_1;
wire na523_1;
wire na525_1;
wire na528_2;
wire na531_1;
wire na533_2;
wire na535_1;
wire na536_1;
wire na538_1;
wire na539_1;
wire na544_1;
wire na545_2;
wire na548_1;
wire na549_1;
wire na551_1;
wire na556_1;
wire na557_2;
wire na560_1;
wire na564_1;
wire na567_1;
wire na568_1;
wire na569_1;
wire na570_1;
wire na571_2;
wire na572_1;
wire na574_1;
wire na578_1;
wire na581_1;
wire na582_1;
wire na583_2;
wire na586_1;
wire na587_1;
wire na590_1;
wire na594_1;
wire na595_1;
wire na596_1;
wire na600_2;
wire na603_1;
wire na604_1;
wire na608_1;
wire na611_1;
wire na612_1;
wire na613_1;
wire na616_1;
wire na617_1;
wire na617_2;
wire na620_1;
wire na625_1;
wire na628_1;
wire na632_1;
wire na635_1;
wire na639_1;
wire na641_1;
wire na642_1;
wire na643_1;
wire na646_1;
wire na648_1;
wire na649_1;
wire na652_1;
wire na655_1;
wire na656_1;
wire na660_1;
wire na662_1;
wire na662_2;
wire na664_1;
wire na665_1;
wire na669_1;
wire na671_1;
wire na672_1;
wire na677_1;
wire na678_1;
wire na683_1;
wire na684_1;
wire na684_2;
wire na687_1;
wire na688_1;
wire na689_1;
wire na693_1;
wire na695_1;
wire na698_1;
wire na702_1;
wire na706_1;
wire na707_1;
wire na708_1;
wire na711_1;
wire na714_1;
wire na718_1;
wire na719_1;
wire na721_1;
wire na726_1;
wire na727_1;
wire na728_1;
wire na731_1;
wire na732_2;
wire na736_1;
wire na737_1;
wire na738_1;
wire na739_1;
wire na740_1;
wire na741_1;
wire na774_1;
wire na775_1;
wire na776_1;
wire na777_1;
wire na778_1;
wire na780_1;
wire na781_1;
wire na782_1;
wire na783_1;
wire na785_1;
wire na787_1;
wire na788_1;
wire na789_1;
wire na790_1;
wire na792_1;
wire na793_1;
wire na794_1;
wire na795_1;
wire na796_1;
wire na797_1;
wire na800_1;
wire na802_1;
wire na803_1;
wire na805_1;
wire na806_1;
wire na809_1;
wire na810_1;
wire na812_1;
wire na813_1;
wire na815_1;
wire na817_1;
wire na819_1;
wire na821_1;
wire na822_1;
wire na824_1;
wire na825_1;
wire na827_1;
wire na828_1;
wire na830_1;
wire na831_1;
wire na833_1;
wire na834_1;
wire na836_1;
wire na838_1;
wire na839_1;
wire na841_1;
wire na843_1;
wire na845_1;
wire na847_1;
wire na848_1;
wire na850_1;
wire na853_1;
wire na853_1_i;
wire na853_2;
wire na853_4;
wire na855_1;
wire na855_1_i;
wire na855_2;
wire na855_4;
wire na857_1;
wire na857_1_i;
wire na857_2;
wire na857_4;
wire na859_1;
wire na859_1_i;
wire na859_2;
wire na859_4;
wire na861_1;
wire na861_1_i;
wire na861_2;
wire na861_4;
wire na862_1;
wire na862_1_i;
wire na862_2;
wire na862_4;
wire na864_1;
wire na864_1_i;
wire na864_2;
wire na864_4;
wire na866_1;
wire na866_1_i;
wire na866_2;
wire na866_4;
wire na868_1;
wire na868_1_i;
wire na868_2;
wire na868_4;
wire na870_1;
wire na870_1_i;
wire na870_2;
wire na870_4;
wire na872_1;
wire na872_1_i;
wire na872_2;
wire na872_4;
wire na875_1;
wire na875_1_i;
wire na876_1;
wire na876_1_i;
wire na876_2;
wire na876_4;
wire na878_1;
wire na878_1_i;
wire na878_2;
wire na878_4;
wire na880_1;
wire na880_1_i;
wire na880_2;
wire na880_4;
wire na882_1;
wire na882_1_i;
wire na882_2;
wire na882_4;
wire na883_1;
wire na883_4;
wire na885_1;
wire na885_2;
wire na885_4;
wire na887_1;
wire na887_2;
wire na887_4;
wire na889_1;
wire na889_2;
wire na889_4;
wire na891_1;
wire na891_2;
wire na891_4;
wire na893_1;
wire na893_2;
wire na893_4;
wire na894_1;
wire na894_4;
wire na896_1;
wire na896_2;
wire na896_4;
wire na898_1;
wire na899_1;
wire na899_4;
wire na900_1;
wire na900_4;
wire na901_1;
wire na901_4;
wire na902_1;
wire na902_2;
wire na902_4;
wire na904_1;
wire na904_2;
wire na904_4;
wire na906_1;
wire na906_2;
wire na906_4;
wire na907_1;
wire na907_4;
wire na909_1;
wire na909_2;
wire na909_4;
wire na911_1;
wire na911_2;
wire na911_4;
wire na913_1;
wire na913_2;
wire na913_4;
wire na915_1;
wire na915_2;
wire na915_4;
wire na917_1;
wire na917_2;
wire na917_4;
wire na918_1;
wire na918_2;
wire na918_4;
wire na920_1;
wire na922_1;
wire na922_2;
wire na922_4;
wire na924_1;
wire na924_2;
wire na924_4;
wire na926_1;
wire na926_2;
wire na926_4;
wire na928_1;
wire na928_2;
wire na928_4;
wire na929_1;
wire na929_4;
wire na930_1;
wire na930_4;
wire na931_1;
wire na931_4;
wire na932_1;
wire na932_4;
wire na933_1;
wire na933_4;
wire na934_1;
wire na934_4;
wire na935_1;
wire na935_4;
wire na936_1;
wire na936_4;
wire na937_1;
wire na937_4;
wire na938_1;
wire na938_4;
wire na939_1;
wire na939_4;
wire na940_1;
wire na940_4;
wire na941_1;
wire na941_4;
wire na942_1;
wire na942_4;
wire na943_1;
wire na944_1;
wire na944_4;
wire na945_1;
wire na945_4;
wire na946_1;
wire na946_2;
wire na946_4;
wire na948_1;
wire na948_2;
wire na948_4;
wire na950_1;
wire na950_2;
wire na950_4;
wire na952_1;
wire na952_2;
wire na952_4;
wire na953_1;
wire na953_2;
wire na953_4;
wire na955_1;
wire na955_2;
wire na955_4;
wire na957_1;
wire na957_2;
wire na957_4;
wire na959_1;
wire na959_2;
wire na959_4;
wire na961_1;
wire na961_2;
wire na961_4;
wire na964_1;
wire na964_2;
wire na964_4;
wire na966_1;
wire na966_2;
wire na966_4;
wire na968_1;
wire na968_2;
wire na968_4;
wire na970_1;
wire na970_2;
wire na970_4;
wire na972_1;
wire na972_2;
wire na972_4;
wire na974_1;
wire na974_2;
wire na974_4;
wire na975_1;
wire na975_2;
wire na978_1;
wire na978_2;
wire na978_4;
wire na980_1;
wire na980_2;
wire na980_4;
wire na982_1;
wire na982_2;
wire na982_4;
wire na984_1;
wire na984_2;
wire na984_4;
wire na985_1;
wire na985_2;
wire na985_4;
wire na987_1;
wire na987_2;
wire na987_4;
wire na989_1;
wire na989_2;
wire na989_4;
wire na991_1;
wire na991_2;
wire na991_4;
wire na993_1;
wire na993_2;
wire na993_4;
wire na996_1;
wire na996_2;
wire na996_4;
wire na998_1;
wire na998_2;
wire na998_4;
wire na1000_1;
wire na1000_2;
wire na1000_4;
wire na1002_1;
wire na1002_2;
wire na1002_4;
wire na1004_1;
wire na1004_2;
wire na1004_4;
wire na1006_1;
wire na1006_2;
wire na1006_4;
wire na1007_1;
wire na1007_2;
wire na1007_4;
wire na1009_1;
wire na1009_4;
wire na1011_1;
wire na1011_2;
wire na1011_4;
wire na1013_1;
wire na1013_2;
wire na1013_4;
wire na1015_1;
wire na1015_2;
wire na1015_4;
wire na1018_1;
wire na1023_1;
wire na1023_1_i;
wire na1023_2;
wire na1023_2_i;
wire na1025_1;
wire na1025_1_i;
wire na1027_2;
wire na1027_2_i;
wire na1029_1;
wire na1029_1_i;
wire na1031_2;
wire na1031_2_i;
wire na1033_2;
wire na1033_2_i;
wire na1035_1;
wire na1035_1_i;
wire na1037_1;
wire na1037_1_i;
wire na1039_1;
wire na1039_1_i;
wire na1041_2;
wire na1041_2_i;
wire na1043_1;
wire na1043_1_i;
wire na1045_2;
wire na1045_2_i;
wire na1047_2;
wire na1047_2_i;
wire na1049_2;
wire na1049_2_i;
wire na1051_1;
wire na1051_1_i;
wire na1053_2;
wire na1053_2_i;
wire na1054_1;
wire na1054_1_i;
wire na1055_1;
wire na1055_1_i;
wire na1055_2;
wire na1055_2_i;
wire na1056_1;
wire na1056_1_i;
wire na1058_1;
wire na1058_1_i;
wire na1058_2;
wire na1058_2_i;
wire na1059_1;
wire na1059_1_i;
wire na1059_2;
wire na1059_2_i;
wire na1060_1;
wire na1060_1_i;
wire na1060_2;
wire na1060_2_i;
wire na1061_1;
wire na1061_1_i;
wire na1061_2;
wire na1061_2_i;
wire na1062_1;
wire na1062_1_i;
wire na1062_2;
wire na1062_2_i;
wire na1063_1;
wire na1063_1_i;
wire na1063_2;
wire na1063_2_i;
wire na1064_1;
wire na1064_1_i;
wire na1065_2;
wire na1065_2_i;
wire na1066_1;
wire na1066_1_i;
wire na1067_2;
wire na1067_2_i;
wire na1068_2;
wire na1068_2_i;
wire na1069_2;
wire na1069_2_i;
wire na1070_1;
wire na1070_1_i;
wire na1077_1;
wire na1077_1_i;
wire na1077_2;
wire na1077_2_i;
wire na1079_1;
wire na1079_1_i;
wire na1079_2;
wire na1079_2_i;
wire na1081_1;
wire na1081_1_i;
wire na1081_2;
wire na1081_2_i;
wire na1108_1;
wire na1141_1;
wire na1142_1;
wire na1143_1;
wire na1144_1;
wire na1145_1;
wire na1146_1;
wire na1147_1;
wire na1148_1;
wire na1149_1;
wire na1150_1;
wire na1151_1;
wire na1152_1;
wire na1153_1;
wire na1154_1;
wire na1155_1;
wire na1156_1;
wire na1157_1;
wire na1158_1;
wire na1159_1;
wire na1160_1;
wire na1161_1;
wire na1162_1;
wire na1163_1;
wire na1164_1;
wire na1165_1;
wire na1166_1;
wire na1167_1;
wire na1168_1;
wire na1169_1;
wire na1170_1;
wire na1171_1;
wire na1172_1;
wire na1173_1;
wire na1175_1;
wire na1212_1;
wire na1213_1;
wire na1213_2;
wire na1213_3;
wire na1213_4;
wire na1213_5;
wire na1213_6;
wire na1213_7;
wire na1213_8;
wire na1213_9;
wire na1215_1;
wire na1215_9;
wire na1216_2;
wire na1217_2;
wire na1218_2;
wire na1219_2;
wire na1220_1;
wire na1221_1;
wire na1221_9;
wire na1222_1;
wire na1222_4;
wire na1223_2;
wire na1224_1;
wire na1225_1;
wire na1226_2;
wire na1227_2;
wire na1228_1;
wire na1228_2;
wire na1229_1;
wire na1230_2;
wire na1231_1;
wire na1232_1;
wire na1232_4;
wire na1233_1;
wire na1233_4;
wire na1234_1;
wire na1234_9;
wire na1235_2;
wire na1236_1;
wire na1237_2;
wire na1238_1;
wire na1238_9;
wire na1239_1;
wire na1239_4;
wire na1240_1;
wire na1241_2;
wire na1242_1;
wire na1242_9;
wire na1243_1;
wire na1244_1;
wire na1245_2;
wire na1246_1;
wire na1246_9;
wire na1247_2;
wire na1248_1;
wire na1249_1;
wire na1249_9;
wire na1250_2;
wire na1251_1;
wire na1251_9;
wire na1252_1;
wire na1253_2;
wire na1254_1;
wire na1254_9;
wire na1255_2;
wire na1256_1;
wire na1257_1;
wire na1257_9;
wire na1258_2;
wire na1259_1;
wire na1259_9;
wire na1260_1;
wire na1261_2;
wire na1262_1;
wire na1262_9;
wire na1263_2;
wire na1264_1;
wire na1265_1;
wire na1265_9;
wire na1266_2;
wire na1267_1;
wire na1267_9;
wire na1268_1;
wire na1269_2;
wire na1270_1;
wire na1270_9;
wire na1271_2;
wire na1272_1;
wire na1273_1;
wire na1273_9;
wire na1274_2;
wire na1275_1;
wire na1275_9;
wire na1276_1;
wire na1277_2;
wire na1277_2_i;
wire na1278_1;
wire na1278_1_i;
wire na1278_9;
wire na1279_2;
wire na1279_2_i;
wire na1280_1;
wire na1281_1;
wire na1281_1_i;
wire na1281_9;
wire na1282_2;
wire na1282_2_i;
wire na1283_1;
wire na1283_1_i;
wire na1283_9;
wire na1284_1;
wire na1285_2;
wire na1285_2_i;
wire na1286_1;
wire na1286_1_i;
wire na1286_9;
wire na1287_2;
wire na1287_2_i;
wire na1288_1;
wire na1289_1;
wire na1289_1_i;
wire na1289_9;
wire na1290_2;
wire na1290_2_i;
wire na1291_1;
wire na1291_1_i;
wire na1291_9;
wire na1292_1;
wire na1293_2;
wire na1293_2_i;
wire na1294_1;
wire na1294_1_i;
wire na1294_9;
wire na1295_2;
wire na1295_2_i;
wire na1296_1;
wire na1297_1;
wire na1297_1_i;
wire na1297_9;
wire na1298_2;
wire na1298_2_i;
wire na1299_1;
wire na1299_1_i;
wire na1299_9;
wire na1300_1;
wire na1301_2;
wire na1301_2_i;
wire na1302_1;
wire na1302_1_i;
wire na1302_9;
wire na1303_2;
wire na1303_2_i;
wire na1304_1;
wire na1305_1;
wire na1305_1_i;
wire na1305_9;
wire na1306_2;
wire na1306_2_i;
wire na1307_1;
wire na1307_1_i;
wire na1307_9;
wire na1308_1;
wire na1309_2;
wire na1309_2_i;
wire na1310_1;
wire na1310_1_i;
wire na1310_9;
wire na1311_2;
wire na1311_2_i;
wire na1312_1;
wire na1313_1;
wire na1313_1_i;
wire na1313_9;
wire na1314_2;
wire na1314_2_i;
wire na1315_1;
wire na1315_1_i;
wire na1315_9;
wire na1316_1;
wire na1317_2;
wire na1317_2_i;
wire na1318_1;
wire na1318_1_i;
wire na1318_9;
wire na1319_2;
wire na1320_1;
wire na1321_1;
wire na1321_9;
wire na1322_2;
wire na1323_1;
wire na1323_9;
wire na1324_2;
wire na1325_1;
wire na1325_9;
wire na1326_1;
wire na1327_1;
wire na1328_2;
wire na1329_1;
wire na1330_1;
wire na1330_9;
wire na1331_1;
wire na1332_1;
wire na1333_1;
wire na1334_1;
wire na1334_9;
wire na1335_2;
wire na1336_1;
wire na1337_1;
wire na1338_2;
wire na1339_1;
wire na1339_9;
wire na1340_2;
wire na1341_1;
wire na1341_2;
wire na1342_1;
wire na1343_1;
wire na1343_9;
wire na1344_2;
wire na1345_1;
wire na1345_9;
wire na1346_2;
wire na1347_1;
wire na1348_1;
wire na1349_1;
wire na1350_1;
wire na1351_1;
wire na1352_1;
wire na1353_1;
wire na1354_2;
wire na1355_1;
wire na1356_1;
wire na1356_2;
wire na1357_2;
wire na1358_1;
wire na1358_9;
wire na1359_1;
wire na1360_2;
wire na1361_2;
wire na1362_2;
wire na1363_1;
wire na1363_9;
wire na1364_1;
wire na1365_1;
wire na1366_1;
wire na1367_2;
wire na1368_1;
wire na1368_9;
wire na1369_2;
wire na1370_1;
wire na1371_1;
wire na1371_9;
wire na1372_1;
wire na1373_2;
wire na1374_1;
wire na1375_2;
wire na1376_1;
wire na1376_2;
wire na1377_1;
wire na1378_1;
wire na1378_9;
wire na1379_2;
wire na1380_2;
wire na1381_1;
wire na1381_9;
wire na1382_1;
wire na1383_1;
wire na1384_1;
wire na1385_2;
wire na1386_1;
wire na1387_1;
wire na1387_9;
wire na1388_2;
wire na1389_1;
wire na1390_1;
wire na1391_2;
wire na1392_1;
wire na1392_9;
wire na1393_1;
wire na1394_2;
wire na1395_2;
wire na1396_1;
wire na1397_1;
wire na1397_2;
wire na1398_2;
wire na1399_1;
wire na1400_1;
wire na1401_1;
wire na1402_1;
wire na1403_1;
wire na1403_9;
wire na1404_2;
wire na1405_1;
wire na1405_9;
wire na1406_2;
wire na1407_2;
wire na1408_2;
wire na1409_1;
wire na1409_9;
wire na1410_1;
wire na1411_2;
wire na1412_1;
wire na1413_1;
wire na1414_1;
wire na1415_1;
wire na1416_2;
wire na1417_1;
wire na1418_1;
wire na1419_1;
wire na1419_9;
wire na1420_1;
wire na1421_1;
wire na1421_2;
wire na1422_2;
wire na1423_2;
wire na1424_1;
wire na1425_1;
wire na1425_9;
wire na1426_2;
wire na1427_1;
wire na1428_1;
wire na1429_1;
wire na1430_2;
wire na1430_2_i;
wire na1431_1;
wire na1432_1;
wire na1433_1;
wire na1433_1_i;
wire na1433_9;
wire na1434_1;
wire na1435_1;
wire na1436_2;
wire na1436_2_i;
wire na1437_1;
wire na1438_2;
wire na1439_2;
wire na1440_1;
wire na1441_1;
wire na1442_1;
wire na1442_1_i;
wire na1442_9;
wire na1443_1;
wire na1444_1;
wire na1445_1;
wire na1446_1;
wire na1447_2;
wire na1447_2_i;
wire na1448_1;
wire na1449_1;
wire na1450_1;
wire na1450_2;
wire na1451_1;
wire na1452_1;
wire na1452_1_i;
wire na1452_9;
wire na1453_2;
wire na1454_2;
wire na1454_2_i;
wire na1455_1;
wire na1455_1_i;
wire na1455_9;
wire na1456_2;
wire na1457_2;
wire na1458_1;
wire na1459_2;
wire na1459_2_i;
wire na1460_1;
wire na1461_1;
wire na1462_1;
wire na1463_1;
wire na1463_1_i;
wire na1463_9;
wire na1464_1;
wire na1465_2;
wire na1466_2;
wire na1467_1;
wire na1468_2;
wire na1468_2_i;
wire na1469_1;
wire na1470_1;
wire na1471_1;
wire na1472_1;
wire na1473_2;
wire na1474_1;
wire na1474_1_i;
wire na1474_9;
wire na1475_2;
wire na1475_2_i;
wire na1476_1;
wire na1477_1;
wire na1478_1;
wire na1478_1_i;
wire na1478_9;
wire na1479_1;
wire na1480_2;
wire na1480_2_i;
wire na1481_1;
wire na1482_1;
wire na1483_1;
wire na1484_1;
wire na1484_1_i;
wire na1484_9;
wire na1485_1;
wire na1486_1;
wire na1487_2;
wire na1488_1;
wire na1489_1;
wire na1490_1;
wire na1491_2;
wire na1491_2_i;
wire na1492_1;
wire na1492_1_i;
wire na1492_9;
wire na1493_2;
wire na1493_2_i;
wire na1494_1;
wire na1495_1;
wire na1496_1;
wire na1496_1_i;
wire na1496_9;
wire na1497_2;
wire na1497_2_i;
wire na1498_1;
wire na1499_1;
wire na1500_2;
wire na1501_1;
wire na1502_1;
wire na1503_1;
wire na1503_1_i;
wire na1503_9;
wire na1504_2;
wire na1504_2_i;
wire na1505_1;
wire na1506_2;
wire na1507_1;
wire na1508_1;
wire na1509_1;
wire na1509_1_i;
wire na1509_9;
wire na1510_2;
wire na1510_2_i;
wire na1511_1;
wire na1512_2;
wire na1513_1;
wire na1514_1;
wire na1514_1_i;
wire na1514_9;
wire na1515_1;
wire na1516_2;
wire na1516_2_i;
wire na1517_1;
wire na1517_1_i;
wire na1517_9;
wire na1518_2;
wire na1518_2_i;
wire na1519_1;
wire na1519_1_i;
wire na1519_9;
wire na1520_2;
wire na1520_2_i;
wire na1521_1;
wire na1522_2;
wire na1523_2;
wire na1524_1;
wire na1525_1;
wire na1525_1_i;
wire na1525_9;
wire na1526_2;
wire na1527_2;
wire na1528_2;
wire na1529_1;
wire na1530_1;
wire na1530_9;
wire na1531_1;
wire na1532_1;
wire na1533_2;
wire na1534_1;
wire na1534_9;
wire na1535_2;
wire na1536_1;
wire na1537_1;
wire na1538_1;
wire na1539_1;
wire na1539_9;
wire na1540_2;
wire na1541_1;
wire na1542_2;
wire na1543_1;
wire na1544_1;
wire na1545_1;
wire na1546_1;
wire na1546_9;
wire na1547_1;
wire na1548_1;
wire na1553_1;
wire na1555_2;
wire na1556_2;
wire na1557_1;
wire na1558_2;
wire na1559_2;
wire na1561_1;
wire na1563_2;
wire na1564_1;
wire na1565_2;
wire na1566_1;
wire na1567_1;
wire na1568_1;
wire na1568_2;
wire na1569_1;
wire na1570_1;
wire na1574_2;
wire na1576_1;
wire na1577_1;
wire na1580_2;
wire na1581_1;
wire na1582_2;
wire na1584_1;
wire na1585_2;
wire na1588_2;
wire na1589_1;
wire na1590_2;
wire na1592_1;
wire na1593_1;
wire na1596_2;
wire na1597_1;
wire na1598_2;
wire na1599_1;
wire na1599_2;
wire na1603_1;
wire na1606_2;
wire na1607_1;
wire na1608_1;
wire na1612_1;
wire na1614_2;
wire na1615_2;
wire na1616_1;
wire na1617_1;
wire na1618_1;
wire na1619_1;
wire na1619_2;
wire na1623_1;
wire na1624_1;
wire na1626_2;
wire na1630_2;
wire na1631_1;
wire na1632_2;
wire na1635_1;
wire na1636_2;
wire na1637_1;
wire na1642_1;
wire na1643_2;
wire na1651_1;
wire na1652_1;
wire na1657_1;
wire na1658_2;
wire na1662_1;
wire na1667_1;
wire na1668_1;
wire na1668_2;
wire na1671_1;
wire na1673_1;
wire na1676_2;
wire na1681_1;
wire na1682_1;
wire na1682_2;
wire na1683_1;
wire na1687_2;
wire na1692_1;
wire na1695_1;
wire na1698_1;
wire na1703_2;
wire na1705_1;
wire na1705_2;
wire na1708_1;
wire na1710_1;
wire na1712_1;
wire na1715_1;
wire na1717_1;
wire na1718_1;
wire na1720_1;
wire na1721_2;
wire na1730_1;
wire na1731_1;
wire na1732_1;
wire na1734_2;
wire na1735_2;
wire na1738_2;
wire na1739_1;
wire na1741_2;
wire na1742_1;
wire na1743_1;
wire na1745_1;
wire na1750_1;
wire na1751_1;
wire na1753_2;
wire na1754_1;
wire na1756_1;
wire na1757_1;
wire na1758_1;
wire na1760_1;
wire na1761_1;
wire na1766_2;
wire na1767_1;
wire na1769_1;
wire na1769_2;
wire na1770_1;
wire na1772_1;
wire na1772_2;
wire na1773_1;
wire na1775_1;
wire na1778_2;
wire na1779_1;
wire na1782_1;
wire na1782_2;
wire na1783_1;
wire na1788_2;
wire na1790_2;
wire na1791_1;
wire na1793_1;
wire na1795_1;
wire na1796_1;
wire na1797_2;
wire na1798_2;
wire na1799_2;
wire na1800_2;
wire na1801_2;
wire na1802_2;
wire na1803_2;
wire na1804_2;
wire na1805_2;
wire na1806_2;
wire na1807_2;
wire na1808_2;
wire na1809_2;
wire na1810_2;
wire na1811_2;
wire na1812_2;
wire na1813_2;
wire na1814_2;
wire na1815_2;
wire na1816_2;
wire na1817_2;
wire na1818_2;
wire na1819_2;
wire na1820_2;
wire na1821_2;
wire na1822_2;
wire na1823_2;
wire na1824_2;
wire na1825_2;
wire na1826_2;
wire na1827_2;
wire na1828_2;
wire na1829_2;
wire na1830_2;
wire na1831_2;
wire na1832_2;
wire na1833_2;
wire na1834_2;
wire na1835_2;
wire na1836_2;
wire na1837_2;
wire na1838_2;
wire na1839_2;
wire na1840_2;
wire na1841_2;
wire na1842_2;
wire na1843_2;
wire na1844_2;
wire na1845_2;
wire na1846_2;
wire na1847_2;
wire na1848_2;
wire na1849_2;
wire na1850_2;
wire na1851_2;
wire na1852_2;
wire na1853_2;
wire na1854_2;
wire na1855_2;
wire na1856_2;
wire na1857_2;
wire na1858_2;
wire na1859_2;
wire na1860_2;
wire na1861_2;
wire na1862_2;
wire na1863_2;
wire na1864_2;
wire na1865_2;
wire na1866_2;
wire na1867_2;
wire na1868_2;
wire na1869_2;
wire na1870_2;
wire na1871_2;
wire na1872_2;
wire na1873_2;
wire na1874_2;
wire na1875_2;
wire na1876_2;
wire na1877_2;
wire na1878_2;
wire na1879_2;
wire na1880_2;
wire na1881_2;
wire na1882_2;
wire na1883_2;
wire na1884_2;
wire na1885_2;
wire na1886_2;
wire na1887_2;
wire na1888_2;
wire na1889_2;
wire na1890_2;
wire na1891_2;
wire na1892_2;
wire na1893_2;
wire na1894_2;
wire na1895_2;
wire na1896_2;
wire na1897_2;
wire na1898_2;
wire na1899_2;
wire na1900_2;
wire na1901_2;
wire na1902_2;
wire na1903_2;
wire na1904_2;
wire na1905_2;
wire na1906_2;
wire na1907_2;
wire na1908_2;
wire na1909_2;
wire na1910_2;
wire na1911_2;
wire na1912_2;
wire na1913_2;
wire na1914_2;
wire na1915_2;
wire na1916_2;
wire na1917_2;
wire na1918_2;
wire na1919_2;
wire na1920_2;
wire na1921_2;
wire na1922_2;
wire na1923_2;
wire na1924_2;
wire na1925_2;
wire na1926_2;
wire na1927_2;
wire na1928_2;
wire na1929_2;
wire na1930_2;
wire na1931_2;
wire na1932_2;
wire na1933_2;
wire na1934_2;
wire na1935_2;
wire na1936_2;
wire na1937_2;
wire na1938_2;
wire na1939_2;
wire na1940_2;
wire na1941_2;
wire na1942_2;
wire na1943_2;
wire na1944_2;
wire na1945_2;
wire na1946_2;
wire na1947_2;
wire na1948_2;
wire na1949_2;
wire na1950_2;
wire na1951_2;
wire na1952_2;
wire na1953_2;
wire na1954_2;
wire na1955_2;
wire na1956_2;
wire na1957_2;
wire na1958_2;
wire na1959_2;
wire na1960_2;
wire na1961_2;
wire na1962_2;
wire na1963_2;
wire na1964_2;
wire na1965_2;
wire na1966_2;
wire na1967_2;
wire na1968_2;
wire na1969_2;
wire na1970_2;
wire na1971_2;
wire na1972_2;
wire na1973_2;
wire na1974_2;
wire na1975_2;
wire na1976_2;
wire na1977_2;
wire na1978_2;
wire na1979_2;
wire na1980_2;
wire na1981_2;
wire na1982_2;
wire na1983_2;
wire na1984_2;
wire na1985_2;
wire na1986_2;
wire na1987_2;
wire na1988_2;
wire na1989_2;
wire na1990_2;
wire na1991_2;
wire na1992_2;
wire na1993_2;
wire na1994_2;
wire na1995_2;
wire na1996_2;
wire na1997_2;
wire na1998_2;
wire na1999_2;
wire na2000_2;
wire na2001_2;
wire na2002_2;
wire na2003_2;
wire na2004_2;
wire na2005_2;
wire na2006_2;
wire na2007_2;
wire na2008_2;
wire na2009_2;
wire na2010_2;
wire na2011_2;
wire na2012_2;
wire na2013_2;
wire na2014_2;
wire na2015_2;
wire na2016_2;
wire na2017_2;
wire na2018_2;
wire na2019_2;
wire na2020_2;
wire na2021_2;
wire na2022_2;
wire na2023_2;
wire na2024_2;
wire na2025_2;
wire na2026_2;
wire na2027_2;
wire na2028_2;
wire na2029_2;
wire na2030_2;
wire na2031_2;
wire na2032_2;
wire na2033_2;
wire na2034_2;
wire na2035_2;
wire na2036_2;
wire na2037_2;
wire na2038_2;
wire na2039_2;
wire na2040_2;
wire na2041_2;
wire na2042_2;
wire na2043_2;
wire na2044_2;
wire na2045_2;
wire na2046_2;
wire na2047_2;
wire na2048_2;
wire na2049_2;
wire na2050_2;
wire na2051_2;
wire na2052_2;
wire na2053_2;
wire na2054_2;
wire na2055_2;
wire na2056_2;
wire na2057_2;
wire na2058_2;
wire na2059_2;
wire na2060_2;
wire na2061_2;
wire na2062_2;
wire na2063_2;
wire na2064_2;
wire na2065_2;
wire na2066_2;
wire na2067_2;
wire na2068_2;
wire na2069_2;
wire na2070_2;
wire na2071_2;
wire na2072_2;
wire na2073_2;
wire na2074_2;
wire na2075_2;
wire na2076_2;
wire na2077_2;
wire na2078_2;
wire na2079_2;
wire na2080_2;
wire na2081_2;
wire na2082_2;
wire na2083_2;
wire na2084_2;
wire na2085_2;
wire na2086_2;
wire na2087_2;
wire na2088_2;
wire na2089_2;
wire na2090_2;
wire na2091_2;
wire na2092_2;
wire na2093_2;
wire na2094_2;
wire na2095_2;
wire na2096_2;
wire na2097_2;
wire na2098_2;
wire na2099_2;
wire na2100_2;
wire na2101_2;
wire na2102_2;
wire na2103_2;
wire na2104_2;
wire na2105_2;
wire na2106_2;
wire na2107_2;
wire na2108_2;
wire na2109_2;
wire na2110_2;
wire na2111_2;
wire na2112_2;
wire na2113_2;
wire na2114_2;
wire na2115_2;
wire na2116_2;
wire mem_rbusy;
wire mem_rstrb;
wire mem_wbusy;
wire na1213_10;
wire na1213_11;
wire na1213_12;
wire na1213_13;
wire na1213_14;
wire na1213_15;
wire na1213_16;
wire na1213_17;
wire na1213_18;
wire na1213_19;
wire na1213_20;
wire na1213_89;
wire na1213_90;
wire na1213_91;
wire na1213_92;
wire na1213_93;
wire na1213_94;
wire na1213_95;
wire na1213_96;
wire na1213_97;
wire na1213_98;
wire na1213_99;
wire na1214_21;
wire na1214_22;
wire na1214_23;
wire na1214_24;
wire na1214_25;
wire na1214_26;
wire na1214_27;
wire na1214_28;
wire na1214_29;
wire na1214_30;
wire na1214_31;
wire na1214_32;
wire na1214_33;
wire na1214_34;
wire na1214_35;
wire na1214_36;
wire na1214_37;
wire na1214_38;
wire na1214_39;
wire na1214_40;
wire na1217_10;
wire na1219_10;
wire na1230_10;
wire na1237_10;
wire na1241_10;
wire na1245_10;
wire na1247_10;
wire na1250_10;
wire na1253_10;
wire na1255_10;
wire na1258_10;
wire na1261_10;
wire na1263_10;
wire na1266_10;
wire na1269_10;
wire na1271_10;
wire na1274_10;
wire na1277_10;
wire na1279_10;
wire na1282_10;
wire na1285_10;
wire na1287_10;
wire na1290_10;
wire na1293_10;
wire na1295_10;
wire na1298_10;
wire na1301_10;
wire na1303_10;
wire na1306_10;
wire na1309_10;
wire na1311_10;
wire na1314_10;
wire na1317_10;
wire na1319_10;
wire na1322_10;
wire na1324_10;
wire na1328_10;
wire na1335_10;
wire na1338_10;
wire na1340_10;
wire na1344_10;
wire na1354_10;
wire na1360_10;
wire na1367_10;
wire na1369_10;
wire na1373_10;
wire na1380_10;
wire na1385_10;
wire na1388_10;
wire na1398_10;
wire na1404_10;
wire na1406_10;
wire na1416_10;
wire na1423_10;
wire na1430_10;
wire na1436_10;
wire na1447_10;
wire na1454_10;
wire na1459_10;
wire na1468_10;
wire na1475_10;
wire na1480_10;
wire na1491_10;
wire na1493_10;
wire na1497_10;
wire na1504_10;
wire na1510_10;
wire na1516_10;
wire na1518_10;
wire na1520_10;
wire na1526_10;
wire na1533_10;
wire na1535_10;
wire na1540_10;
wire na1797_10;
wire na1798_10;
wire na1799_10;
wire na1800_10;
wire na1801_10;
wire na1802_10;
wire na1803_10;
wire na1804_10;
wire na1805_10;
wire na1806_10;
wire na1807_10;
wire na1808_10;
wire na1809_10;
wire na1810_10;
wire na1811_10;
wire na1812_10;
wire na1813_10;
wire na1814_10;
wire na1815_10;
wire na1816_10;
wire na1817_10;
wire na1818_10;
wire na1819_10;
wire na1820_10;
wire na1821_10;
wire na1822_10;
wire na1823_10;
wire na1824_10;
wire na1825_10;
wire na1826_10;
wire na1827_10;
wire na1828_10;
wire na1829_10;
wire na1830_10;
wire na1831_10;
wire na1832_10;
wire na1833_10;
wire na1834_10;
wire na1835_10;
wire na1836_10;
wire na1837_10;
wire na1838_10;
wire na1839_10;
wire na1840_10;
wire na1841_10;
wire na1842_10;
wire na1843_10;
wire na1844_10;
wire na1845_10;
wire na1846_10;
wire na1847_10;
wire na1848_10;
wire na1849_10;
wire na1850_10;
wire na1851_10;
wire na1852_10;
wire na1853_10;
wire na1854_10;
wire na1855_10;
wire na1856_10;
wire na1857_10;
wire na1858_10;
wire na1859_10;
wire na1860_10;
wire na1861_10;
wire na1862_10;
wire na1863_10;
wire na1864_10;
wire na1865_10;
wire na1213_100;
wire na1214_109;
wire na1214_110;
wire na1214_111;
wire na1214_112;
wire na1214_113;
wire na1214_114;
wire na1214_115;
wire na1214_116;
wire na1214_117;
wire na1214_118;
wire na1214_119;
wire na1214_120;

// C_///AND/      x94y67     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1_4 ( .OUT(na1_2), .IN1(1'b1), .IN2(na1212_1), .IN3(~na240_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y63     80'h00_0018_00_0000_0C88_ECFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a2_1 ( .OUT(na2_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na1212_1), .IN7(na1866_2), .IN8(na1216_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x85y71     80'h00_0060_00_0000_0C08_FFCE
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3_4 ( .OUT(na3_2), .IN1(na1141_1), .IN2(na1175_1), .IN3(1'b0), .IN4(na241_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y72     80'h00_0018_00_0040_0A55_0080
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4_1 ( .OUT(na4_1), .IN1(1'b0), .IN2(1'b0), .IN3(na6_1), .IN4(na5_1), .IN5(~na1058_2), .IN6(1'b0), .IN7(~na1302_1), .IN8(1'b0),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x86y68     80'h00_0078_00_0000_0C88_C1A3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5_1 ( .OUT(na5_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1053_2), .IN6(~na1054_1), .IN7(1'b1), .IN8(na1056_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5_4 ( .OUT(na5_2), .IN1(1'b1), .IN2(~na1054_1), .IN3(na1055_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x82y67     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6_1 ( .OUT(na6_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2019_2), .IN6(1'b0), .IN7(na1055_2), .IN8(1'b0),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y68     80'h00_0018_00_0040_0A55_0080
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7_1 ( .OUT(na7_1), .IN1(1'b0), .IN2(1'b0), .IN3(na6_1), .IN4(na5_1), .IN5(~na1059_2), .IN6(1'b0), .IN7(~na1301_2), .IN8(1'b0),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y68     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1), .IN1(1'b1), .IN2(na9_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1060_2), .IN8(~na1299_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x71y62     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9_4 ( .OUT(na9_2), .IN1(1'b1), .IN2(1'b1), .IN3(na6_1), .IN4(na5_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                   .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y67     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a10_1 ( .OUT(na10_1), .IN1(1'b1), .IN2(na9_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2027_2), .IN8(~na1298_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y64     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a11_1 ( .OUT(na11_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1874_2), .IN5(~na1062_2), .IN6(1'b0), .IN7(~na1297_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x75y58     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1295_2), .IN4(~na2041_2), .IN5(1'b1), .IN6(~na9_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y64     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1), .IN1(1'b1), .IN2(na9_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2039_2), .IN8(~na1294_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y59     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a14_1 ( .OUT(na14_1), .IN1(1'b1), .IN2(na9_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2043_2), .IN8(~na1293_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y66     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a15_1 ( .OUT(na15_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1874_2), .IN5(~na1079_1), .IN6(1'b0), .IN7(~na1291_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y66     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a16_1 ( .OUT(na16_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1874_2), .IN5(~na1081_2), .IN6(1'b0), .IN7(~na1290_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x71y66     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a17_1 ( .OUT(na17_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na2044_2), .IN4(~na1289_1), .IN5(1'b1), .IN6(na9_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y62     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a18_1 ( .OUT(na18_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na1287_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x77y71     80'h00_0018_00_0040_0C33_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a19_1 ( .OUT(na19_1), .IN1(~na2056_2), .IN2(~na1063_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na9_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y68     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a20_1 ( .OUT(na20_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na2055_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y67     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a21_1 ( .OUT(na21_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na1283_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y67     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na1282_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y61     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a23_1 ( .OUT(na23_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na2051_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x68y64     80'h00_0018_00_0040_0C33_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a24_1 ( .OUT(na24_1), .IN1(~na2050_2), .IN2(~na1063_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na9_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y70     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a25_1 ( .OUT(na25_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na1278_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x73y70     80'h00_0018_00_0040_0C33_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a26_1 ( .OUT(na26_1), .IN1(~na2047_2), .IN2(~na1063_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na9_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y67     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na2072_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x68y66     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a28_1 ( .OUT(na28_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na2070_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x63y65     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a29_1 ( .OUT(na29_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na1315_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x63y66     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a30_1 ( .OUT(na30_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na1314_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x74y70     80'h00_0018_00_0040_0C33_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a31_1 ( .OUT(na31_1), .IN1(~na2066_2), .IN2(~na1063_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na9_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x63y67     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a32_1 ( .OUT(na32_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na2065_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x63y68     80'h00_0018_00_0040_0C33_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_1 ( .OUT(na33_1), .IN1(~na2064_2), .IN2(~na1063_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na9_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x69y73     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a34_1 ( .OUT(na34_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na1309_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y73     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a35_1 ( .OUT(na35_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na2063_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y72     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na2062_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y70     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a37_1 ( .OUT(na37_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1874_2), .IN5(1'b0), .IN6(~na1063_2), .IN7(1'b0), .IN8(~na1305_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x79y71     80'h00_0018_00_0040_0CAA_8F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a38_1 ( .OUT(na38_1), .IN1(1'b0), .IN2(~na1063_2), .IN3(1'b0), .IN4(~na1303_2), .IN5(1'b1), .IN6(1'b1), .IN7(na6_1), .IN8(na5_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x77y62     80'h00_0018_00_0000_0888_BFE5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_1 ( .OUT(na39_1), .IN1(~na1220_1), .IN2(1'b0), .IN3(na240_2), .IN4(na241_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1055_1),
                    .IN8(~na5_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a40 ( .PCLK0(na40_1), .PCLK1(_d0), .PCLK2(_d1), .PCLK3(_d2), .CLK0(na1108_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0), .SER_CLK(1'b0),
                  .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_ORAND/D///      x92y69     80'h00_FE00_00_0000_0C88_CDFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a42_1 ( .OUT(na42_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na46_1), .IN6(na1228_2), .IN7(1'b0), .IN8(na1212_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a42_2 ( .OUT(na42_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na42_1_i) );
// C_AND///AND/      x84y70     80'h00_0078_00_0000_0C88_54C3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a44_1 ( .OUT(na44_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1053_2), .IN6(na1902_2), .IN7(~na1055_2),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a44_4 ( .OUT(na44_2), .IN1(1'b1), .IN2(~na1054_1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y67     80'h00_0018_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1054_1), .IN7(~na1055_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y61     80'h00_0018_00_0040_0A55_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a46_1 ( .OUT(na46_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na42_1), .IN4(1'b1), .IN5(~na1141_1), .IN6(1'b0), .IN7(~na1218_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x77y69     80'h00_F600_80_0000_0C08_FF38
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a47_4 ( .OUT(na47_2_i), .IN1(na47_2), .IN2(na1212_1), .IN3(1'b1), .IN4(~na44_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a47_5 ( .OUT(na47_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na47_2_i) );
// C_AND///AND/      x86y64     80'h00_0078_00_0000_0C88_8285
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a49_1 ( .OUT(na49_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1053_2), .IN6(~na2020_2), .IN7(na1055_2), .IN8(na1056_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a49_4 ( .OUT(na49_2), .IN1(~na2019_2), .IN2(1'b1), .IN3(na1055_2), .IN4(na5_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x88y72     80'h00_F600_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a50_1 ( .OUT(na50_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1212_1), .IN7(1'b1), .IN8(na241_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a50_2 ( .OUT(na50_1), .CLK(na1018_1), .EN(~na2_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na50_1_i) );
// C_MX2a////      x82y79     80'h00_0018_00_0040_0C45_1000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1), .IN1(na47_2), .IN2(1'b0), .IN3(~na76_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na42_1), .IN8(~na50_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x82y75     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a76_1 ( .OUT(na76_1), .IN1(1'b1), .IN2(na1228_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na883_1), .IN8(~na2046_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x84y81     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a77_1 ( .OUT(na77_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na1913_2), .IN7(~na1229_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x81y69     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na44_2), .IN5(1'b0), .IN6(~na952_2), .IN7(1'b0), .IN8(~na79_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y64     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a79_1 ( .OUT(na79_1), .IN1(~na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1912_2), .IN6(na929_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x91y67     80'h00_0018_00_0040_0C8A_3F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1), .IN1(1'b0), .IN2(na1231_1), .IN3(1'b0), .IN4(~na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na49_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x92y82     80'h00_0018_00_0040_0A55_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a81_1 ( .OUT(na81_1), .IN1(na84_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1243_1), .IN5(~na85_1), .IN6(1'b0), .IN7(~na1905_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x80y69     80'h00_0060_00_0000_0C08_FFC1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a83_4 ( .OUT(na83_2), .IN1(~na1064_1), .IN2(~na1063_1), .IN3(1'b1), .IN4(na1065_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x73y63     80'h00_0078_00_0000_0C88_C8A3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a84_1 ( .OUT(na84_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1064_1), .IN6(na1063_1), .IN7(1'b1), .IN8(na1065_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a84_4 ( .OUT(na84_2), .IN1(1'b1), .IN2(~na349_1), .IN3(na83_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x71y61     80'h00_0018_00_0000_0C88_C2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a85_1 ( .OUT(na85_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(1'b1), .IN8(na1065_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x91y62     80'h00_0018_00_0040_0AAA_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a86_1 ( .OUT(na86_1), .IN1(1'b1), .IN2(~na101_2), .IN3(na90_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na101_1), .IN7(1'b0), .IN8(~na102_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x79y64     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1064_1), .IN6(na1063_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x68y63     80'h00_0018_00_0000_0888_8888
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1), .IN1(na99_1), .IN2(na92_1), .IN3(na97_1), .IN4(na100_1), .IN5(na99_2), .IN6(na92_2), .IN7(na97_2),
                    .IN8(na100_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x67y62     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a92_1 ( .OUT(na92_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2008_2), .IN6(~na2009_2), .IN7(~na998_2),
                    .IN8(~na996_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a92_4 ( .OUT(na92_2), .IN1(~na2006_2), .IN2(~na2007_2), .IN3(~na993_2), .IN4(~na991_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x72y61     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a97_1 ( .OUT(na97_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2015_2), .IN6(~na2016_2), .IN7(~na1013_2),
                    .IN8(~na1011_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a97_4 ( .OUT(na97_2), .IN1(~na2012_2), .IN2(~na2014_2), .IN3(~na1007_2), .IN4(~na1004_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x67y65     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a99_1 ( .OUT(na99_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2004_2), .IN6(~na2005_2), .IN7(~na989_2),
                    .IN8(~na987_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a99_4 ( .OUT(na99_2), .IN1(~na2010_2), .IN2(~na2011_2), .IN3(~na1002_2), .IN4(~na1000_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x72y60     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a100_1 ( .OUT(na100_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2017_2), .IN6(~na2003_2), .IN7(~na985_2),
                     .IN8(~na1015_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a100_4 ( .OUT(na100_2), .IN1(~na2002_2), .IN2(~na2013_2), .IN3(~na1006_2), .IN4(~na984_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x79y66     80'h00_0078_00_0000_0C88_34CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a101_1 ( .OUT(na101_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1064_1), .IN6(na1063_1), .IN7(1'b1), .IN8(~na1065_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a101_4 ( .OUT(na101_2), .IN1(1'b1), .IN2(na349_1), .IN3(1'b1), .IN4(na102_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x80y70     80'h00_0078_00_0000_0C88_31CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a102_1 ( .OUT(na102_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1064_1), .IN6(~na1063_1), .IN7(1'b1), .IN8(~na1065_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a102_4 ( .OUT(na102_2), .IN1(1'b1), .IN2(na89_1), .IN3(1'b1), .IN4(na1065_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x94y82     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a106_1 ( .OUT(na106_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na1916_2), .IN7(1'b0), .IN8(~na1236_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x87y71     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a107_1 ( .OUT(na107_1), .IN1(1'b1), .IN2(~na1899_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na974_1), .IN6(~na108_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y60     80'h00_0018_00_0040_0A32_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a108_1 ( .OUT(na108_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na940_1), .IN6(~na1916_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x100y81     80'h00_0060_00_0000_0C08_FF3B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a111_4 ( .OUT(na111_2), .IN1(na1235_2), .IN2(~na249_1), .IN3(1'b0), .IN4(~na1240_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y65     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a112_1 ( .OUT(na112_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na44_2), .IN5(~na974_2), .IN6(1'b0), .IN7(~na113_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y63     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a113_1 ( .OUT(na113_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na2001_2), .IN6(na918_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x100y55     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a116_1 ( .OUT(na116_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na1915_2), .IN7(1'b0), .IN8(~na1244_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x87y63     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a117_1 ( .OUT(na117_1), .IN1(1'b1), .IN2(na1899_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na118_1), .IN6(~na978_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y57     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a118_1 ( .OUT(na118_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na945_1), .IN6(na918_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x100y59     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a121_4 ( .OUT(na121_2), .IN1(na1235_2), .IN2(~na252_2), .IN3(~na1248_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y61     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a122_1 ( .OUT(na122_1), .IN1(1'b1), .IN2(na1899_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na123_1), .IN6(~na978_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y69     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a123_1 ( .OUT(na123_1), .IN1(~na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na922_1), .IN6(na946_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x100y57     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a126_1 ( .OUT(na126_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na252_1), .IN7(~na1252_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y59     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a127_1 ( .OUT(na127_1), .IN1(1'b1), .IN2(~na1899_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na980_1), .IN6(~na128_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y68     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1), .IN1(~na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na922_2), .IN6(na946_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x98y59     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a131_4 ( .OUT(na131_2), .IN1(na1235_2), .IN2(~na254_2), .IN3(~na1256_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y69     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a132_1 ( .OUT(na132_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na44_2), .IN5(~na980_2), .IN6(1'b0), .IN7(~na133_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y67     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a133_1 ( .OUT(na133_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na948_1), .IN6(na924_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x100y59     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a136_1 ( .OUT(na136_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na254_1), .IN7(1'b0), .IN8(~na1260_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x91y73     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a137_1 ( .OUT(na137_1), .IN1(1'b1), .IN2(na1899_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na138_1), .IN6(~na982_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y65     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na948_2), .IN6(na924_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x100y63     80'h00_0060_00_0000_0C08_FF3B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a141_4 ( .OUT(na141_2), .IN1(na1235_2), .IN2(~na256_2), .IN3(1'b0), .IN4(~na1264_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y73     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a142_1 ( .OUT(na142_1), .IN1(1'b1), .IN2(na1899_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na143_1), .IN6(~na982_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y69     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a143_1 ( .OUT(na143_1), .IN1(~na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na926_1), .IN6(na950_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y76     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a146_1 ( .OUT(na146_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na256_1), .IN7(1'b0), .IN8(~na1268_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x87y69     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a147_1 ( .OUT(na147_1), .IN1(1'b1), .IN2(~na1899_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na953_1), .IN6(~na148_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y58     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a148_1 ( .OUT(na148_1), .IN1(~na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na926_2), .IN6(na950_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x84y81     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a151_4 ( .OUT(na151_2), .IN1(na1235_2), .IN2(~na258_2), .IN3(~na1272_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y67     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a152_1 ( .OUT(na152_1), .IN1(1'b1), .IN2(~na1899_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na953_2), .IN6(~na153_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x97y66     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a153_1 ( .OUT(na153_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na930_1), .IN6(na928_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x90y82     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a156_1 ( .OUT(na156_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na258_1), .IN7(~na1276_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y73     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a157_1 ( .OUT(na157_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na44_2), .IN5(1'b0), .IN6(~na955_1), .IN7(1'b0), .IN8(~na158_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y70     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a158_1 ( .OUT(na158_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1998_2), .IN6(na928_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x86y81     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a161_4 ( .OUT(na161_2), .IN1(na1235_2), .IN2(~na1920_2), .IN3(~na1280_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x81y75     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a162_1 ( .OUT(na162_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na44_2), .IN5(1'b0), .IN6(~na955_2), .IN7(1'b0), .IN8(~na163_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y70     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a163_1 ( .OUT(na163_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na932_1), .IN6(na1995_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x75y54     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a166_1 ( .OUT(na166_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na1919_2), .IN7(~na1284_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y77     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a167_1 ( .OUT(na167_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na44_2), .IN5(~na957_1), .IN6(1'b0), .IN7(~na168_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x86y69     80'h00_0018_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a168_1 ( .OUT(na168_1), .IN1(na909_2), .IN2(na933_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na80_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x93y80     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a171_1 ( .OUT(na171_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na262_2), .IN7(~na1288_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y75     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a172_1 ( .OUT(na172_1), .IN1(1'b1), .IN2(~na1899_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na957_2), .IN6(~na173_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x91y72     80'h00_0018_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a173_1 ( .OUT(na173_1), .IN1(na934_1), .IN2(na911_1), .IN3(1'b0), .IN4(1'b0), .IN5(na80_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y81     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a176_1 ( .OUT(na176_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na262_1), .IN7(1'b0), .IN8(~na1292_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y77     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a177_1 ( .OUT(na177_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na44_2), .IN5(1'b0), .IN6(~na959_1), .IN7(1'b0), .IN8(~na178_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x94y70     80'h00_0018_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a178_1 ( .OUT(na178_1), .IN1(na1999_2), .IN2(na911_2), .IN3(1'b0), .IN4(1'b0), .IN5(na80_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x87y82     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a181_4 ( .OUT(na181_2), .IN1(na1235_2), .IN2(~na264_2), .IN3(~na1296_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y75     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_1 ( .OUT(na182_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na44_2), .IN5(1'b0), .IN6(~na959_2), .IN7(1'b0), .IN8(~na183_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y72     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a183_1 ( .OUT(na183_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na936_1), .IN6(na1996_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x82y82     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a186_1 ( .OUT(na186_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na264_1), .IN7(1'b0), .IN8(~na1300_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x91y75     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a187_1 ( .OUT(na187_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na44_2), .IN5(~na961_1), .IN6(1'b0), .IN7(~na188_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x94y71     80'h00_0018_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a188_1 ( .OUT(na188_1), .IN1(na913_2), .IN2(na937_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na80_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x89y81     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a191_4 ( .OUT(na191_2), .IN1(na1235_2), .IN2(~na266_2), .IN3(~na1304_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x91y77     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a192_1 ( .OUT(na192_1), .IN1(1'b1), .IN2(~na1899_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na961_2), .IN6(~na193_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x91y74     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a193_1 ( .OUT(na193_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na938_1), .IN6(na915_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x99y81     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a196_1 ( .OUT(na196_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na266_1), .IN7(~na1308_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x87y79     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a197_1 ( .OUT(na197_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na44_2), .IN5(1'b0), .IN6(~na964_1), .IN7(1'b0), .IN8(~na198_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x94y72     80'h00_0018_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a198_1 ( .OUT(na198_1), .IN1(na2000_2), .IN2(na915_2), .IN3(1'b0), .IN4(1'b0), .IN5(na80_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x98y81     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a201_4 ( .OUT(na201_2), .IN1(na1235_2), .IN2(~na268_2), .IN3(~na1312_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x93y77     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a202_1 ( .OUT(na202_1), .IN1(1'b1), .IN2(na1899_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na203_1), .IN6(~na964_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x95y75     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a203_1 ( .OUT(na203_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na941_1), .IN6(na1997_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x100y81     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a206_1 ( .OUT(na206_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1235_2), .IN6(~na268_1), .IN7(1'b0), .IN8(~na1316_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y79     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a207_1 ( .OUT(na207_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na44_2), .IN5(~na966_1), .IN6(1'b0), .IN7(~na208_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x96y75     80'h00_0018_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a208_1 ( .OUT(na208_1), .IN1(na917_2), .IN2(na942_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na80_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x99y81     80'h00_0060_00_0000_0C08_FF3B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a211_4 ( .OUT(na211_2), .IN1(na1235_2), .IN2(~na269_2), .IN3(1'b0), .IN4(~na1320_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y77     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a212_1 ( .OUT(na212_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na44_2), .IN5(~na966_2), .IN6(1'b0), .IN7(~na213_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x96y71     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a213_1 ( .OUT(na213_1), .IN1(na80_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na943_1), .IN6(na920_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y61     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a216_1 ( .OUT(na216_1), .IN1(1'b1), .IN2(~na1970_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1302_1), .IN8(na2061_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x63y63     80'h00_0018_00_0040_0C05_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a217_1 ( .OUT(na217_1), .IN1(na2060_2), .IN2(1'b0), .IN3(na1301_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na883_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y46     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a218_1 ( .OUT(na218_1), .IN1(1'b1), .IN2(na1970_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2059_2), .IN8(na1299_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x77y46     80'h00_0018_00_0040_0C0A_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a219_1 ( .OUT(na219_1), .IN1(1'b0), .IN2(na2058_2), .IN3(1'b0), .IN4(na1298_2), .IN5(1'b1), .IN6(1'b1), .IN7(na883_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y47     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a220_1 ( .OUT(na220_1), .IN1(1'b1), .IN2(~na1970_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1297_1), .IN8(na2057_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x79y45     80'h00_0018_00_0040_0C05_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a221_1 ( .OUT(na221_1), .IN1(na2054_2), .IN2(1'b0), .IN3(na1295_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na883_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y46     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a222_1 ( .OUT(na222_1), .IN1(1'b1), .IN2(na1970_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2053_2), .IN8(na1294_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x79y48     80'h00_0018_00_0040_0C0A_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a223_1 ( .OUT(na223_1), .IN1(1'b0), .IN2(na2052_2), .IN3(1'b0), .IN4(na1293_2), .IN5(1'b1), .IN6(1'b1), .IN7(na883_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y46     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a224_1 ( .OUT(na224_1), .IN1(1'b1), .IN2(~na1982_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1302_1), .IN8(na2051_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x86y46     80'h00_0018_00_0040_0C05_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a225_1 ( .OUT(na225_1), .IN1(na2050_2), .IN2(1'b0), .IN3(na1301_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y45     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a226_1 ( .OUT(na226_1), .IN1(1'b1), .IN2(na1982_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2049_2), .IN8(na1299_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x66y51     80'h00_0018_00_0040_0C0A_CF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a227_1 ( .OUT(na227_1), .IN1(1'b0), .IN2(na2048_2), .IN3(1'b0), .IN4(na1298_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x66y47     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a228_1 ( .OUT(na228_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na894_1), .IN5(na2071_2), .IN6(1'b0), .IN7(na1297_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x66y52     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a229_1 ( .OUT(na229_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na894_1), .IN5(na2069_2), .IN6(1'b0), .IN7(na1295_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x68y53     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a230_1 ( .OUT(na230_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na894_1), .IN5(1'b0), .IN6(na2068_2), .IN7(1'b0), .IN8(na1294_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x66y54     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a231_1 ( .OUT(na231_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na894_1), .IN5(1'b0), .IN6(na2067_2), .IN7(1'b0), .IN8(na1293_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x67y55     80'h00_0018_00_0040_0C05_1000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a232_1 ( .OUT(na232_1), .IN1(na216_1), .IN2(1'b0), .IN3(na1313_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na883_1), .IN8(~na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x66y56     80'h00_0018_00_0040_0C05_1000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a233_1 ( .OUT(na233_1), .IN1(na217_1), .IN2(1'b0), .IN3(na1311_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na883_1), .IN8(~na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x67y54     80'h00_0018_00_0040_0C0A_1F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a234_1 ( .OUT(na234_1), .IN1(1'b0), .IN2(na218_1), .IN3(1'b0), .IN4(na1310_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na883_1), .IN8(~na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x65y53     80'h00_0018_00_0040_0C0A_1F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a235_1 ( .OUT(na235_1), .IN1(1'b0), .IN2(na219_1), .IN3(1'b0), .IN4(na1309_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na883_1), .IN8(~na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x66y53     80'h00_0018_00_0040_0C05_1000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a236_1 ( .OUT(na236_1), .IN1(na220_1), .IN2(1'b0), .IN3(na1307_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na883_1), .IN8(~na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x65y55     80'h00_0018_00_0040_0C05_1000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a237_1 ( .OUT(na237_1), .IN1(na221_1), .IN2(1'b0), .IN3(na1306_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na883_1), .IN8(~na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x65y59     80'h00_0018_00_0040_0C0A_1F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a238_1 ( .OUT(na238_1), .IN1(1'b0), .IN2(na222_1), .IN3(1'b0), .IN4(na1305_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na883_1), .IN8(~na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x65y58     80'h00_0018_00_0040_0C0A_1F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a239_1 ( .OUT(na239_1), .IN1(1'b0), .IN2(na223_1), .IN3(1'b0), .IN4(na1303_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na883_1), .IN8(~na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x82y65     80'h00_FE18_00_0000_0888_AFF4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a240_1 ( .OUT(na240_1), .IN1(~na1141_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na42_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a240_5 ( .OUT(na240_2), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na240_1) );
// C_ORAND*/D///      x82y68     80'h00_FE00_00_0000_0788_FC75
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a241_1 ( .OUT(na241_1_i), .IN1(~na3_2), .IN2(1'b0), .IN3(~na240_2), .IN4(~na44_1), .IN5(1'b0), .IN6(na1212_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a241_2 ( .OUT(na241_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na241_1_i) );
// C_///AND/D      x88y65     80'h00_F600_80_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a247_4 ( .OUT(na247_2_i), .IN1(~na78_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a247_5 ( .OUT(na247_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na247_2_i) );
// C_AND/D///      x97y70     80'h00_F600_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a249_1 ( .OUT(na249_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na112_1), .IN6(na1212_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a249_2 ( .OUT(na249_1), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na249_1_i) );
// C_AND/D//AND/D      x90y64     80'h00_F600_80_0000_0C88_F4F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a250_1 ( .OUT(na250_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na117_1), .IN6(na1212_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a250_2 ( .OUT(na250_1), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na250_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a250_4 ( .OUT(na250_2_i), .IN1(~na107_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a250_5 ( .OUT(na250_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na250_2_i) );
// C_AND/D//AND/D      x97y62     80'h00_F600_80_0000_0C88_F4F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a252_1 ( .OUT(na252_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na127_1), .IN6(na1212_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a252_2 ( .OUT(na252_1), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na252_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a252_4 ( .OUT(na252_2_i), .IN1(~na122_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a252_5 ( .OUT(na252_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na252_2_i) );
// C_AND/D//AND/D      x97y64     80'h00_F600_80_0000_0C88_F4F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a254_1 ( .OUT(na254_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na137_1), .IN6(na1212_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a254_2 ( .OUT(na254_1), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na254_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a254_4 ( .OUT(na254_2_i), .IN1(~na132_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a254_5 ( .OUT(na254_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na254_2_i) );
// C_AND/D//AND/D      x91y70     80'h00_F600_80_0000_0C88_F4F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a256_1 ( .OUT(na256_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na147_1), .IN6(na1212_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a256_2 ( .OUT(na256_1), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na256_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a256_4 ( .OUT(na256_2_i), .IN1(~na142_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a256_5 ( .OUT(na256_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na256_2_i) );
// C_AND/D//AND/D      x89y76     80'h00_F600_80_0000_0C88_F4F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a258_1 ( .OUT(na258_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na157_1), .IN6(na1212_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a258_2 ( .OUT(na258_1), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na258_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a258_4 ( .OUT(na258_2_i), .IN1(~na152_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a258_5 ( .OUT(na258_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na258_2_i) );
// C_AND/D//AND/D      x90y76     80'h00_F600_80_0000_0C88_F4F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a260_1 ( .OUT(na260_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na167_1), .IN6(na1212_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a260_2 ( .OUT(na260_1), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na260_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a260_4 ( .OUT(na260_2_i), .IN1(~na162_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a260_5 ( .OUT(na260_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na260_2_i) );
// C_AND/D//AND/D      x93y76     80'h00_F600_80_0000_0C88_F4F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a262_1 ( .OUT(na262_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na177_1), .IN6(na1212_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a262_2 ( .OUT(na262_1), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na262_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a262_4 ( .OUT(na262_2_i), .IN1(~na172_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a262_5 ( .OUT(na262_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na262_2_i) );
// C_AND/D//AND/D      x89y78     80'h00_F600_80_0000_0C88_F4F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a264_1 ( .OUT(na264_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na187_1), .IN6(na1212_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a264_2 ( .OUT(na264_1), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na264_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a264_4 ( .OUT(na264_2_i), .IN1(~na182_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a264_5 ( .OUT(na264_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na264_2_i) );
// C_AND/D//AND/D      x91y78     80'h00_F600_80_0000_0C88_F4F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a266_1 ( .OUT(na266_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na197_1), .IN6(na1212_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a266_2 ( .OUT(na266_1), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na266_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a266_4 ( .OUT(na266_2_i), .IN1(~na192_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a266_5 ( .OUT(na266_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na266_2_i) );
// C_AND/D//AND/D      x93y78     80'h00_F600_80_0000_0C88_F4F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a268_1 ( .OUT(na268_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na207_1), .IN6(na1212_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a268_2 ( .OUT(na268_1), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na268_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a268_4 ( .OUT(na268_2_i), .IN1(~na202_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a268_5 ( .OUT(na268_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na268_2_i) );
// C_///AND/D      x95y78     80'h00_F600_80_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a269_4 ( .OUT(na269_2_i), .IN1(~na212_1), .IN2(na1212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a269_5 ( .OUT(na269_2), .CLK(na1018_1), .EN(~na1_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na269_2_i) );
// C_ORAND////      x79y63     80'h00_0018_00_0000_0888_7DBD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a270_1 ( .OUT(na270_1), .IN1(~na47_2), .IN2(na2075_2), .IN3(na1326_1), .IN4(~na350_1), .IN5(~na1341_2), .IN6(na1342_1), .IN7(~na2018_2),
                     .IN8(~na350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x68y67     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a272_1 ( .OUT(na272_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1496_1), .IN8(~na1497_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x63y69     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a273_1 ( .OUT(na273_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1493_2), .IN8(~na1503_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y69     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a274_1 ( .OUT(na274_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1504_2), .IN8(~na1492_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y70     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a275_1 ( .OUT(na275_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1509_1), .IN8(~na1491_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y74     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a276_1 ( .OUT(na276_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na277_1), .IN6(na280_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y65     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a277_1 ( .OUT(na277_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na278_1), .IN6(na279_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x61y69     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a278_1 ( .OUT(na278_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1484_1), .IN8(~na1510_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y74     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a279_1 ( .OUT(na279_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1480_2), .IN8(~na1514_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y68     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a280_1 ( .OUT(na280_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na281_1), .IN6(na282_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y65     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a281_1 ( .OUT(na281_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1516_2), .IN8(~na1478_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x63y72     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a282_1 ( .OUT(na282_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1517_1), .IN8(~na1475_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y72     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a283_1 ( .OUT(na283_1), .IN1(1'b1), .IN2(na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(na291_1), .IN6(na1931_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x81y65     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_1 ( .OUT(na284_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na285_1), .IN6(na288_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y71     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a285_1 ( .OUT(na285_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na286_1), .IN6(na287_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x63y61     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a286_1 ( .OUT(na286_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1474_1), .IN8(~na1518_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y66     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a287_1 ( .OUT(na287_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1468_2), .IN8(~na1519_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x69y74     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a288_1 ( .OUT(na288_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na289_1), .IN6(na290_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y67     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a289_1 ( .OUT(na289_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1520_2), .IN8(~na1463_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y68     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a290_1 ( .OUT(na290_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1525_1), .IN8(~na1459_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y65     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a291_1 ( .OUT(na291_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na292_1), .IN6(na295_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y73     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a292_1 ( .OUT(na292_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na293_1), .IN6(na294_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y69     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a293_1 ( .OUT(na293_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1455_1), .IN8(~na1430_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y70     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a294_1 ( .OUT(na294_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1454_2), .IN8(~na1433_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y76     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a295_1 ( .OUT(na295_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na296_1), .IN6(na297_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y73     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a296_1 ( .OUT(na296_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1436_2), .IN8(~na1452_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y74     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a297_1 ( .OUT(na297_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1442_1), .IN8(~na1447_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x82y72     80'h00_0018_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a298_1 ( .OUT(na298_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na314_2), .IN6(na299_2), .IN7(1'b0), .IN8(~na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y66     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a299_4 ( .OUT(na299_2), .IN1(1'b1), .IN2(1'b1), .IN3(na10_1), .IN4(~na516_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y76     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a300_1 ( .OUT(na300_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na7_1), .IN5(1'b0), .IN6(na304_1), .IN7(1'b0), .IN8(na301_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x68y72     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a301_1 ( .OUT(na301_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na302_1), .IN6(na1933_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y73     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a302_1 ( .OUT(na302_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1442_1), .IN8(~na1447_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y76     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a303_1 ( .OUT(na303_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1436_2), .IN8(~na1452_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y76     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a304_1 ( .OUT(na304_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1868_2), .IN5(na306_1), .IN6(1'b0), .IN7(na305_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x64y73     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a305_1 ( .OUT(na305_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1454_2), .IN8(~na1433_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x63y73     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a306_1 ( .OUT(na306_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1455_1), .IN4(~na1430_2), .IN5(1'b1), .IN6(~na101_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y74     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a307_1 ( .OUT(na307_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na308_1), .IN6(na1935_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x77y73     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a308_1 ( .OUT(na308_1), .IN1(na310_1), .IN2(na309_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na4_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x65y62     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a309_1 ( .OUT(na309_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1525_1), .IN8(~na1459_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y77     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a310_1 ( .OUT(na310_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1520_2), .IN8(~na1463_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y75     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a311_1 ( .OUT(na311_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1868_2), .IN5(1'b0), .IN6(na312_1), .IN7(1'b0), .IN8(na313_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x69y78     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a312_1 ( .OUT(na312_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1468_2), .IN8(~na1519_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x70y76     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a313_1 ( .OUT(na313_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1474_1), .IN4(~na1518_2), .IN5(1'b1), .IN6(~na101_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x87y67     80'h00_0060_00_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a314_4 ( .OUT(na314_2), .IN1(na315_2), .IN2(na322_1), .IN3(~na10_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x77y67     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a315_4 ( .OUT(na315_2), .IN1(1'b1), .IN2(na8_1), .IN3(na1332_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y73     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a316_1 ( .OUT(na316_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na317_1), .IN8(na318_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y77     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a317_1 ( .OUT(na317_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1517_1), .IN8(~na1475_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y78     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a318_1 ( .OUT(na318_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1516_2), .IN8(~na1478_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x72y76     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a319_1 ( .OUT(na319_1), .IN1(1'b0), .IN2(1'b0), .IN3(na320_1), .IN4(na321_1), .IN5(1'b1), .IN6(~na4_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y75     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a320_1 ( .OUT(na320_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1480_2), .IN8(~na1514_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y78     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a321_1 ( .OUT(na321_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1484_1), .IN8(~na1510_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x79y62     80'h00_0018_00_0000_0C88_E3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a322_1 ( .OUT(na322_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na8_1), .IN7(na326_1), .IN8(na323_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x78y78     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a323_1 ( .OUT(na323_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na406_1), .IN8(na7_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y75     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a324_1 ( .OUT(na324_1), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1509_1), .IN8(~na1491_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x70y74     80'h00_0018_00_0040_0CCC_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a325_1 ( .OUT(na325_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1504_2), .IN4(~na1492_1), .IN5(1'b1), .IN6(na101_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y61     80'h00_0018_00_0040_0ACC_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a326_1 ( .OUT(na326_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b1), .IN4(~na7_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na328_1), .IN8(~na1939_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y67     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a327_1 ( .OUT(na327_1), .IN1(1'b1), .IN2(~na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1496_1), .IN8(~na1497_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x72y65     80'h00_0018_00_0040_0CCC_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a328_1 ( .OUT(na328_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1493_2), .IN4(~na1503_1), .IN5(1'b1), .IN6(~na101_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x82y70     80'h00_0018_00_0040_0A51_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a330_1 ( .OUT(na330_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na11_1), .IN5(~na333_2), .IN6(1'b0), .IN7(na331_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x86y65     80'h00_0018_00_0040_0C15_8000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a331_1 ( .OUT(na331_1), .IN1(~na333_2), .IN2(1'b0), .IN3(na332_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na10_1), .IN8(na1873_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x80y71     80'h00_0018_00_0040_0C15_8000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a332_1 ( .OUT(na332_1), .IN1(~na333_2), .IN2(1'b0), .IN3(na327_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1867_2), .IN8(na7_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x85y73     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a333_4 ( .OUT(na333_2), .IN1(na1081_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1497_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x79y61     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a334_1 ( .OUT(na334_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1336_1), .IN7(1'b1), .IN8(na102_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x74y62     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a335_1 ( .OUT(na335_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1081_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1056_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x74y61     80'h00_0018_00_0040_0A76_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a336_1 ( .OUT(na336_1), .IN1(1'b1), .IN2(~na2106_2), .IN3(1'b1), .IN4(na1868_2), .IN5(na85_1), .IN6(~na2074_2), .IN7(~na1337_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y58     80'h00_0018_00_0040_0AC0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a342_1 ( .OUT(na342_1), .IN1(1'b1), .IN2(na1982_2), .IN3(1'b1), .IN4(na343_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1142_1), .IN8(na1150_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x80y62     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a343_1 ( .OUT(na343_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1064_1), .IN6(1'b0), .IN7(~na883_1), .IN8(na2030_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x76y60     80'h00_0018_00_0040_0C55_3000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a344_1 ( .OUT(na344_1), .IN1(~na1159_1), .IN2(1'b0), .IN3(~na1172_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x84y61     80'h00_0018_00_0000_0C88_18FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a346_1 ( .OUT(na346_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1053_2), .IN6(na1870_2), .IN7(~na1055_2),
                     .IN8(~na1056_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x84y58     80'h00_0078_00_0000_0C88_123C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a348_1 ( .OUT(na348_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1064_1), .IN6(~na349_1), .IN7(~na2029_2),
                     .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a348_4 ( .OUT(na348_2), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(~na330_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x63y74     80'h00_0018_00_0040_0CB9_3500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a349_1 ( .OUT(na349_1), .IN1(~na2107_2), .IN2(1'b1), .IN3(1'b0), .IN4(~na1497_2), .IN5(~na38_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na1243_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x82y62     80'h00_0078_00_0000_0C88_458A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a350_1 ( .OUT(na350_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1053_2), .IN6(1'b1), .IN7(~na1055_2), .IN8(na5_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a350_4 ( .OUT(na350_2), .IN1(na2019_2), .IN2(1'b1), .IN3(na1055_2), .IN4(na5_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x74y59     80'h00_0018_00_0000_0EEE_5CDA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a351_1 ( .OUT(na351_1), .IN1(na1357_2), .IN2(1'b0), .IN3(~na1356_1), .IN4(na1361_2), .IN5(1'b0), .IN6(na1346_2), .IN7(~na1356_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y70     80'h00_0018_00_0000_0888_CFB5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a352_1 ( .OUT(na352_1), .IN1(~na364_1), .IN2(1'b0), .IN3(na1734_2), .IN4(~na11_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0), .IN8(na102_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y68     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a353_1 ( .OUT(na353_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na281_1), .IN6(na279_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y72     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a354_1 ( .OUT(na354_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na286_1), .IN6(na282_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x69y75     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a355_1 ( .OUT(na355_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na274_1), .IN6(~na1930_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y68     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a356_1 ( .OUT(na356_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na278_1), .IN6(na275_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x83y80     80'h00_0018_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a357_1 ( .OUT(na357_1), .IN1(1'b1), .IN2(na8_1), .IN3(~na10_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na361_1), .IN8(na358_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y80     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a358_1 ( .OUT(na358_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na359_1), .IN6(na360_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y71     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a359_1 ( .OUT(na359_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na289_1), .IN6(na287_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y72     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a360_1 ( .OUT(na360_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na293_1), .IN6(na290_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y81     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a361_1 ( .OUT(na361_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na362_1), .IN6(na363_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x71y77     80'h00_0018_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a362_1 ( .OUT(na362_1), .IN1(na296_1), .IN2(na294_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na4_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y80     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a363_1 ( .OUT(na363_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na302_1), .IN6(na297_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x91y79     80'h00_0018_00_0000_0888_3FDE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a364_1 ( .OUT(na364_1), .IN1(na1875_2), .IN2(na1350_1), .IN3(~na10_1), .IN4(na1348_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(~na11_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y80     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a367_1 ( .OUT(na367_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na305_1), .IN8(na303_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y79     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a368_1 ( .OUT(na368_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na306_1), .IN6(na309_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x76y81     80'h00_0018_00_0040_0ACC_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a369_1 ( .OUT(na369_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b1), .IN4(~na1873_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na371_1),
                     .IN8(~na1948_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y72     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a370_1 ( .OUT(na370_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na310_1), .IN6(na312_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x74y71     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a371_1 ( .OUT(na371_1), .IN1(1'b0), .IN2(1'b0), .IN3(na317_1), .IN4(na313_1), .IN5(1'b1), .IN6(na4_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y74     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a374_1 ( .OUT(na374_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na320_1), .IN8(na318_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x76y73     80'h00_0018_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a375_1 ( .OUT(na375_1), .IN1(1'b0), .IN2(1'b0), .IN3(na324_1), .IN4(na321_1), .IN5(1'b1), .IN6(na4_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x72y69     80'h00_0060_00_0000_0C08_FFE3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a376_4 ( .OUT(na376_2), .IN1(1'b0), .IN2(~na8_1), .IN3(na1949_2), .IN4(na377_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x80y64     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a377_4 ( .OUT(na377_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1353_1), .IN4(na7_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x83y63     80'h00_0018_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a378_1 ( .OUT(na378_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b1), .IN4(na7_1), .IN5(na333_2), .IN6(~na1938_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x83y69     80'h00_0018_00_0040_0C15_8000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a380_1 ( .OUT(na380_1), .IN1(~na333_2), .IN2(1'b0), .IN3(na381_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na10_1), .IN8(na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x88y73     80'h00_0018_00_0040_0C15_8000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a381_1 ( .OUT(na381_1), .IN1(~na333_2), .IN2(1'b0), .IN3(na382_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1872_2), .IN8(na7_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y65     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a382_1 ( .OUT(na382_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na328_1), .IN8(na1939_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x81y60     80'h00_0018_00_0000_0888_F773
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a386_1 ( .OUT(na386_1), .IN1(1'b0), .IN2(~na388_1), .IN3(~na510_2), .IN4(~na1359_1), .IN5(~na1064_1), .IN6(~na1143_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y58     80'h00_0018_00_0040_0AC0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a388_1 ( .OUT(na388_1), .IN1(na1981_2), .IN2(1'b1), .IN3(1'b1), .IN4(na343_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1143_1), .IN8(na1151_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x83y70     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a390_1 ( .OUT(na390_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na399_1), .IN6(na391_2), .IN7(1'b0), .IN8(na102_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x83y70     80'h00_0060_00_0000_0C08_FFCE
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a391_4 ( .OUT(na391_2), .IN1(na392_1), .IN2(na1364_1), .IN3(1'b0), .IN4(na11_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y81     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a392_1 ( .OUT(na392_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na10_1), .IN8(na1365_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y71     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a393_1 ( .OUT(na393_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na7_1), .IN5(na277_1), .IN6(1'b0), .IN7(na394_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x68y65     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a394_1 ( .OUT(na394_1), .IN1(1'b1), .IN2(~na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(na274_1), .IN6(na275_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y75     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a395_1 ( .OUT(na395_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na285_1), .IN6(na280_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y76     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a396_1 ( .OUT(na396_1), .IN1(1'b1), .IN2(na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(na398_1), .IN6(na397_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y76     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a397_1 ( .OUT(na397_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na292_1), .IN6(na288_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y81     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a398_1 ( .OUT(na398_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na7_1), .IN5(1'b0), .IN6(na295_1), .IN7(1'b0), .IN8(na301_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x95y79     80'h00_0018_00_0000_0C88_3EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a399_1 ( .OUT(na399_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na400_1), .IN6(na403_1), .IN7(1'b0), .IN8(~na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y81     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a400_1 ( .OUT(na400_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na10_1), .IN8(~na538_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y82     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a401_1 ( .OUT(na401_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na308_1), .IN6(na304_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x78y82     80'h00_0018_00_0040_0C05_3000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a402_1 ( .OUT(na402_1), .IN1(na311_1), .IN2(1'b0), .IN3(na316_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na7_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y80     80'h00_0018_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a403_1 ( .OUT(na403_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1876_2), .IN7(~na470_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y77     80'h00_0018_00_0040_0A51_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a404_1 ( .OUT(na404_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na7_1), .IN5(~na333_2), .IN6(1'b0), .IN7(na382_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x78y73     80'h00_0018_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a406_1 ( .OUT(na406_1), .IN1(1'b0), .IN2(1'b0), .IN3(na324_1), .IN4(na325_1), .IN5(1'b1), .IN6(~na4_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x68y61     80'h00_0060_00_0000_0C08_FFEC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a407_4 ( .OUT(na407_2), .IN1(1'b0), .IN2(na101_1), .IN3(na1372_1), .IN4(na410_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y72     80'h00_0018_00_0040_0A51_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a408_1 ( .OUT(na408_1), .IN1(1'b0), .IN2(1'b0), .IN3(na10_1), .IN4(1'b1), .IN5(~na333_2), .IN6(1'b0), .IN7(na409_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y79     80'h00_0018_00_0040_0A51_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a409_1 ( .OUT(na409_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1873_2), .IN5(~na333_2), .IN6(1'b0), .IN7(na1352_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x82y76     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a410_4 ( .OUT(na410_2), .IN1(na333_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na11_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x74y56     80'h00_0018_00_0040_0AC0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a415_1 ( .OUT(na415_1), .IN1(na1981_2), .IN2(1'b1), .IN3(1'b1), .IN4(na343_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1154_1), .IN8(na1152_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y58     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a417_1 ( .OUT(na417_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na894_1), .IN5(~na1161_1), .IN6(1'b0), .IN7(~na1144_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y72     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a418_1 ( .OUT(na418_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na11_1), .IN5(1'b0), .IN6(na425_1), .IN7(1'b0), .IN8(na1382_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y80     80'h00_0018_00_0040_0A33_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a419_1 ( .OUT(na419_1), .IN1(1'b1), .IN2(~na8_1), .IN3(na10_1), .IN4(1'b1), .IN5(~na420_1), .IN6(~na421_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y81     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a420_1 ( .OUT(na420_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na362_1), .IN6(na360_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y82     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a421_1 ( .OUT(na421_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1947_2), .IN6(na367_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x82y66     80'h00_0018_00_0040_0C0A_CF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a423_1 ( .OUT(na423_1), .IN1(1'b0), .IN2(na353_1), .IN3(1'b0), .IN4(na1944_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na7_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x71y78     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a424_1 ( .OUT(na424_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na7_1), .IN5(1'b0), .IN6(na1945_2), .IN7(1'b0), .IN8(na354_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x89y80     80'h00_0018_00_0040_0C05_5000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a425_1 ( .OUT(na425_1), .IN1(na1384_1), .IN2(1'b0), .IN3(na428_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na10_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x86y76     80'h00_0018_00_0040_0ACC_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a427_1 ( .OUT(na427_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b1), .IN4(~na1873_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na371_1),
                     .IN8(~na374_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y83     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a428_1 ( .OUT(na428_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1873_2), .IN5(na1386_1), .IN6(1'b0), .IN7(na332_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x66y75     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a429_4 ( .OUT(na429_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na375_1), .IN4(na7_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y72     80'h00_0018_00_0040_0ACC_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a430_1 ( .OUT(na430_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b1), .IN4(~na7_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na328_1), .IN8(~na325_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x85y67     80'h00_0018_00_0040_0C15_8000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a431_1 ( .OUT(na431_1), .IN1(~na333_2), .IN2(1'b0), .IN3(na432_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na10_1), .IN8(na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y75     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a432_1 ( .OUT(na432_1), .IN1(1'b1), .IN2(na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na333_2), .IN6(na1333_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x74y58     80'h00_0018_00_0000_0888_F773
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a436_1 ( .OUT(na436_1), .IN1(1'b0), .IN2(~na438_1), .IN3(~na510_2), .IN4(~na1393_1), .IN5(~na1064_1), .IN6(~na1165_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x85y60     80'h00_0018_00_0040_0AC0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a438_1 ( .OUT(na438_1), .IN1(na1981_2), .IN2(1'b1), .IN3(1'b1), .IN4(na343_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1165_1), .IN8(na1153_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x82y61     80'h00_0018_00_0000_0EEE_3EAA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a440_1 ( .OUT(na440_1), .IN1(na1412_1), .IN2(1'b0), .IN3(na1407_2), .IN4(1'b0), .IN5(na1408_2), .IN6(na1396_1), .IN7(1'b0),
                     .IN8(~na1411_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x71y55     80'h00_0018_00_0000_0888_1F51
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a441_1 ( .OUT(na441_1), .IN1(~na452_1), .IN2(~na451_1), .IN3(~na1397_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1397_2),
                     .IN8(~na442_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x80y68     80'h00_0018_00_0000_0C88_ECFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a442_1 ( .OUT(na442_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na101_1), .IN7(na1399_1), .IN8(na410_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y81     80'h00_0018_00_0040_0A51_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a443_1 ( .OUT(na443_1), .IN1(1'b0), .IN2(1'b0), .IN3(na10_1), .IN4(1'b1), .IN5(~na333_2), .IN6(1'b0), .IN7(na428_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y69     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a444_1 ( .OUT(na444_1), .IN1(1'b1), .IN2(~na1877_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1400_1), .IN8(na447_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y84     80'h00_0018_00_0040_0A33_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a446_1 ( .OUT(na446_1), .IN1(1'b1), .IN2(~na8_1), .IN3(na10_1), .IN4(1'b1), .IN5(~na291_1), .IN6(~na300_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y74     80'h00_0018_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a447_1 ( .OUT(na447_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na10_1), .IN4(1'b1), .IN5(na1402_1), .IN6(1'b0), .IN7(na432_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x76y78     80'h00_0018_00_0040_0ACC_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a449_1 ( .OUT(na449_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b1), .IN4(~na1873_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na316_1),
                     .IN8(~na319_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x73y52     80'h00_0018_00_0040_0A76_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a451_1 ( .OUT(na451_1), .IN1(1'b1), .IN2(na1877_2), .IN3(~na1484_1), .IN4(1'b1), .IN5(na85_1), .IN6(~na2074_2), .IN7(~na1337_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x81y63     80'h00_0018_00_0000_0C88_2AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a452_1 ( .OUT(na452_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na84_1), .IN6(1'b1), .IN7(na1484_1), .IN8(~na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x71y60     80'h00_0018_00_0040_0CAA_CF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a453_1 ( .OUT(na453_1), .IN1(1'b0), .IN2(~na978_1), .IN3(1'b0), .IN4(~na1011_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na335_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x84y64     80'h00_0018_00_0000_0888_F773
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a456_1 ( .OUT(na456_1), .IN1(1'b0), .IN2(~na458_1), .IN3(~na510_2), .IN4(~na1410_1), .IN5(~na1064_1), .IN6(~na1168_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y56     80'h00_0018_00_0040_0AC0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a458_1 ( .OUT(na458_1), .IN1(na1981_2), .IN2(1'b1), .IN3(1'b1), .IN4(na343_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1168_1), .IN8(na1155_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x90y69     80'h00_0018_00_0040_0C55_3000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a460_1 ( .OUT(na460_1), .IN1(~na1413_1), .IN2(1'b0), .IN3(~na466_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x76y69     80'h00_0018_00_0040_0C0A_3F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a462_1 ( .OUT(na462_1), .IN1(1'b0), .IN2(na353_1), .IN3(1'b0), .IN4(na354_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na7_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x85y78     80'h00_0060_00_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a463_4 ( .OUT(na463_2), .IN1(na464_2), .IN2(na465_1), .IN3(~na10_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x83y79     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a464_4 ( .OUT(na464_2), .IN1(1'b1), .IN2(na8_1), .IN3(~na361_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y80     80'h00_0018_00_0040_0A33_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a465_1 ( .OUT(na465_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b1), .IN4(na1873_2), .IN5(~na368_1), .IN6(~na367_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y75     80'h00_0018_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a466_1 ( .OUT(na466_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na10_1), .IN4(1'b1), .IN5(na1417_1), .IN6(1'b0), .IN7(na409_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x85y77     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a467_4 ( .OUT(na467_2), .IN1(1'b1), .IN2(na8_1), .IN3(na1418_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y80     80'h00_0018_00_0040_0ACC_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a468_1 ( .OUT(na468_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b1), .IN4(~na1873_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na375_1),
                     .IN8(~na374_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x81y71     80'h00_0018_00_0040_0C15_8000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a469_1 ( .OUT(na469_1), .IN1(~na333_2), .IN2(1'b0), .IN3(na470_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na10_1), .IN8(na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x84y77     80'h00_0018_00_0000_0C88_7EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a470_1 ( .OUT(na470_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na404_1), .IN6(na8_1), .IN7(~na1370_1), .IN8(~na1873_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x71y56     80'h00_0018_00_0000_0888_F775
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a474_1 ( .OUT(na474_1), .IN1(~na476_1), .IN2(1'b0), .IN3(~na510_2), .IN4(~na1424_1), .IN5(~na1064_1), .IN6(~na1169_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x75y57     80'h00_0018_00_0040_0A30_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a476_1 ( .OUT(na476_1), .IN1(~na1981_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na343_1), .IN5(na1156_1), .IN6(na1169_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x90y67     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a479_1 ( .OUT(na479_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na11_1), .IN5(~na1427_1), .IN6(1'b0), .IN7(~na482_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y79     80'h00_0018_00_0040_0A33_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a480_1 ( .OUT(na480_1), .IN1(1'b1), .IN2(~na8_1), .IN3(na10_1), .IN4(1'b1), .IN5(~na398_1), .IN6(~na401_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x90y73     80'h00_0018_00_0040_0C05_5000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a482_1 ( .OUT(na482_1), .IN1(na1429_1), .IN2(1'b0), .IN3(na381_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na10_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x76y79     80'h00_0018_00_0040_0ACC_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a484_1 ( .OUT(na484_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b1), .IN4(~na1873_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na406_1),
                     .IN8(~na319_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x89y64     80'h00_0018_00_0000_0C88_ECFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a485_1 ( .OUT(na485_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na101_1), .IN7(na1432_1), .IN8(na410_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x92y75     80'h00_0018_00_0040_0C15_A000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a486_1 ( .OUT(na486_1), .IN1(~na333_2), .IN2(1'b0), .IN3(na2077_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na10_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x73y58     80'h00_0018_00_0000_0888_F775
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a489_1 ( .OUT(na489_1), .IN1(~na491_1), .IN2(1'b0), .IN3(~na510_2), .IN4(~na1437_1), .IN5(~na1064_1), .IN6(~na1170_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x73y57     80'h00_0018_00_0040_0AC0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a491_1 ( .OUT(na491_1), .IN1(na1981_2), .IN2(1'b1), .IN3(1'b1), .IN4(na343_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1170_1), .IN8(na1157_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x84y63     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a493_1 ( .OUT(na493_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na922_2), .IN6(1'b1), .IN7(1'b1), .IN8(na49_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x83y68     80'h00_0060_00_0000_0C08_FFEC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a494_4 ( .OUT(na494_2), .IN1(1'b0), .IN2(na101_1), .IN3(na1441_1), .IN4(na410_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y75     80'h00_0018_00_0040_0A51_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a495_1 ( .OUT(na495_1), .IN1(1'b0), .IN2(1'b0), .IN3(na10_1), .IN4(1'b1), .IN5(~na333_2), .IN6(1'b0), .IN7(na1331_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y67     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a496_1 ( .OUT(na496_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na11_1), .IN5(1'b0), .IN6(na500_1), .IN7(1'b0), .IN8(na1443_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x83y81     80'h00_0018_00_0040_0A33_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a498_1 ( .OUT(na498_1), .IN1(1'b1), .IN2(na8_1), .IN3(na10_1), .IN4(1'b1), .IN5(~na499_1), .IN6(~na421_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y79     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a499_1 ( .OUT(na499_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na368_1), .IN6(na370_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x89y74     80'h00_0018_00_0040_0C0A_AF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a500_1 ( .OUT(na500_1), .IN1(1'b0), .IN2(na501_1), .IN3(1'b0), .IN4(na1445_1), .IN5(1'b1), .IN6(1'b1), .IN7(na10_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x85y82     80'h00_0018_00_0040_0A51_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a501_1 ( .OUT(na501_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1873_2), .IN5(~na333_2), .IN6(1'b0), .IN7(na332_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y80     80'h00_0018_00_0000_0C88_E3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a503_1 ( .OUT(na503_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na8_1), .IN7(na429_2), .IN8(na1953_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x82y49     80'h00_0018_00_0000_0C88_DDFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a508_1 ( .OUT(na508_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1960_2), .IN6(na509_1), .IN7(~na510_2), .IN8(na511_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x79y60     80'h00_0018_00_0040_0C55_3000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a509_1 ( .OUT(na509_1), .IN1(~na1158_1), .IN2(1'b0), .IN3(~na1171_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x68y59     80'h00_0078_00_0000_0C88_51A1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a510_1 ( .OUT(na510_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1064_1), .IN6(~na1063_1), .IN7(~na883_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a510_4 ( .OUT(na510_2), .IN1(~na1064_1), .IN2(~na1063_1), .IN3(na883_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x80y58     80'h00_0018_00_0040_0CAA_CF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a511_1 ( .OUT(na511_1), .IN1(1'b0), .IN2(~na1149_1), .IN3(1'b0), .IN4(~na1167_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na894_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x89y48     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a512_1 ( .OUT(na512_1), .IN1(na1064_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1456_2), .IN6(~na1171_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x85y53     80'h00_0018_00_0000_0EEE_0DEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a513_1 ( .OUT(na513_1), .IN1(1'b0), .IN2(na1461_1), .IN3(na1462_1), .IN4(na1465_2), .IN5(~na1464_1), .IN6(na1457_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x87y70     80'h00_0018_00_0000_0888_DF7C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a514_1 ( .OUT(na514_1), .IN1(1'b0), .IN2(na1911_2), .IN3(~na1460_1), .IN4(~na11_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na495_1),
                     .IN8(na11_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y80     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a516_1 ( .OUT(na516_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1873_2), .IN5(1'b0), .IN6(na300_1), .IN7(1'b0), .IN8(na307_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x91y61     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a517_1 ( .OUT(na517_1), .IN1(1'b1), .IN2(na1877_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na333_2), .IN6(na500_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y55     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a518_1 ( .OUT(na518_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(~na982_1), .IN7(1'b0), .IN8(~na1015_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y45     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a521_1 ( .OUT(na521_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na508_1), .IN8(na102_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y48     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a523_1 ( .OUT(na523_1), .IN1(na1064_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1466_2), .IN6(~na1172_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x86y67     80'h00_0018_00_0040_0C05_3000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a525_1 ( .OUT(na525_1), .IN1(na1467_1), .IN2(1'b0), .IN3(na486_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x81y67     80'h00_0060_00_0000_0C08_FFEC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a528_4 ( .OUT(na528_2), .IN1(1'b0), .IN2(na101_1), .IN3(na1471_1), .IN4(na410_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x96y47     80'h00_0018_00_0000_0888_F757
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a531_1 ( .OUT(na531_1), .IN1(~na2078_2), .IN2(~na89_1), .IN3(~na521_1), .IN4(1'b0), .IN5(~na1064_1), .IN6(~na1173_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y66     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a533_4 ( .OUT(na533_2), .IN1(1'b1), .IN2(na950_1), .IN3(na346_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x90y71     80'h00_0018_00_0000_0888_DF7C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a535_1 ( .OUT(na535_1), .IN1(1'b0), .IN2(na1911_2), .IN3(~na1479_1), .IN4(~na11_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na536_1),
                     .IN8(na11_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x92y73     80'h00_0018_00_0040_0A51_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a536_1 ( .OUT(na536_1), .IN1(1'b0), .IN2(1'b0), .IN3(na10_1), .IN4(1'b1), .IN5(~na333_2), .IN6(1'b0), .IN7(na470_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y80     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a538_1 ( .OUT(na538_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1873_2), .IN5(1'b0), .IN6(na401_1), .IN7(1'b0), .IN8(na402_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x81y67     80'h00_0018_00_0000_0C88_ECFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a539_1 ( .OUT(na539_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na101_1), .IN7(na2099_2), .IN8(na410_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x94y48     80'h00_0018_00_0040_0C33_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a544_1 ( .OUT(na544_1), .IN1(~na1488_1), .IN2(~na1144_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1064_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x83y64     80'h00_0060_00_0000_0C08_FF43
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a545_4 ( .OUT(na545_2), .IN1(1'b1), .IN2(~na548_1), .IN3(~na1489_1), .IN4(na102_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x87y72     80'h00_0018_00_0040_0A51_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a548_1 ( .OUT(na548_1), .IN1(1'b1), .IN2(na1877_2), .IN3(na10_1), .IN4(1'b1), .IN5(~na333_2), .IN6(1'b0), .IN7(na428_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x82y63     80'h00_0018_00_0000_0C88_ECFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a549_1 ( .OUT(na549_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na101_1), .IN7(na2105_2), .IN8(na410_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x96y45     80'h00_0018_00_0000_0888_F757
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a551_1 ( .OUT(na551_1), .IN1(~na2080_2), .IN2(~na89_1), .IN3(~na521_1), .IN4(1'b0), .IN5(~na1064_1), .IN6(~na1145_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y69     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a556_1 ( .OUT(na556_1), .IN1(1'b1), .IN2(na1877_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na333_2), .IN6(na425_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x84y67     80'h00_0060_00_0000_0C08_FF43
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a557_4 ( .OUT(na557_2), .IN1(1'b1), .IN2(~na560_1), .IN3(~na1501_1), .IN4(na102_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x85y72     80'h00_0018_00_0040_0A51_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a560_1 ( .OUT(na560_1), .IN1(1'b1), .IN2(na1877_2), .IN3(na10_1), .IN4(1'b1), .IN5(~na333_2), .IN6(1'b0), .IN7(na432_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x94y47     80'h00_0018_00_0000_0888_F757
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a564_1 ( .OUT(na564_1), .IN1(~na2082_2), .IN2(~na89_1), .IN3(~na521_1), .IN4(1'b0), .IN5(~na1064_1), .IN6(~na1146_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x85y62     80'h00_0018_00_0000_0C88_48FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a567_1 ( .OUT(na567_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1053_2), .IN6(na1870_2), .IN7(~na1055_2),
                     .IN8(na1056_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x87y55     80'h00_0018_00_0000_0EEE_E0DB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a568_1 ( .OUT(na568_1), .IN1(na1524_1), .IN2(~na1523_2), .IN3(~na1527_2), .IN4(na1528_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1522_2),
                     .IN8(na1513_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x87y68     80'h00_0018_00_0000_0888_7B75
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a569_1 ( .OUT(na569_1), .IN1(~na570_1), .IN2(1'b0), .IN3(~na1521_1), .IN4(~na102_1), .IN5(na1965_2), .IN6(~na101_1), .IN7(~na813_1),
                     .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y69     80'h00_0018_00_0000_0C88_45FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a570_1 ( .OUT(na570_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1515_1), .IN6(1'b1), .IN7(~na572_1), .IN8(na102_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x83y76     80'h00_0060_00_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a571_4 ( .OUT(na571_2), .IN1(na467_2), .IN2(na468_1), .IN3(~na10_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x88y71     80'h00_0018_00_0040_0A51_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a572_1 ( .OUT(na572_1), .IN1(1'b1), .IN2(na1877_2), .IN3(na10_1), .IN4(1'b1), .IN5(~na333_2), .IN6(1'b0), .IN7(na409_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x90y65     80'h00_0018_00_0000_0C88_B3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a574_1 ( .OUT(na574_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1952_2), .IN7(na1366_1), .IN8(~na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x95y48     80'h00_0018_00_0000_0888_F757
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a578_1 ( .OUT(na578_1), .IN1(~na2084_2), .IN2(~na89_1), .IN3(~na521_1), .IN4(1'b0), .IN5(~na1064_1), .IN6(~na1147_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x90y61     80'h00_0018_00_0000_0EEE_CBAB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a581_1 ( .OUT(na581_1), .IN1(na1542_2), .IN2(~na1543_1), .IN3(na1544_1), .IN4(1'b0), .IN5(na1538_1), .IN6(~na1541_1), .IN7(1'b0),
                     .IN8(na1529_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x87y66     80'h00_0018_00_0000_0888_7B73
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a582_1 ( .OUT(na582_1), .IN1(1'b0), .IN2(~na583_2), .IN3(~na1537_1), .IN4(~na102_1), .IN5(na587_1), .IN6(~na101_1), .IN7(~na815_1),
                     .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x83y72     80'h00_0060_00_0000_0C08_FF34
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a583_4 ( .OUT(na583_2), .IN1(~na1531_1), .IN2(na1911_2), .IN3(1'b1), .IN4(~na586_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x84y72     80'h00_0018_00_0040_0A51_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a586_1 ( .OUT(na586_1), .IN1(1'b1), .IN2(na1877_2), .IN3(na10_1), .IN4(1'b1), .IN5(~na333_2), .IN6(1'b0), .IN7(na381_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x89y71     80'h00_0018_00_0000_0C88_B3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a587_1 ( .OUT(na587_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1952_2), .IN7(na1536_1), .IN8(~na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x93y47     80'h00_0018_00_0000_0888_F757
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a590_1 ( .OUT(na590_1), .IN1(~na2088_2), .IN2(~na89_1), .IN3(~na521_1), .IN4(1'b0), .IN5(~na1064_1), .IN6(~na1148_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x89y56     80'h00_0018_00_0000_0EEE_EB0D
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a594_1 ( .OUT(na594_1), .IN1(~na1558_2), .IN2(na603_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1557_1), .IN6(~na1556_2), .IN7(na1559_2),
                     .IN8(na1545_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x75y53     80'h00_0018_00_0000_0888_7B73
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a595_1 ( .OUT(na595_1), .IN1(1'b0), .IN2(~na596_1), .IN3(~na1553_1), .IN4(~na102_1), .IN5(na1966_2), .IN6(~na101_1), .IN7(~na817_1),
                     .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x89y70     80'h00_0018_00_0000_0888_F5DC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a596_1 ( .OUT(na596_1), .IN1(1'b0), .IN2(na1911_2), .IN3(~na331_1), .IN4(na11_1), .IN5(~na1547_1), .IN6(1'b0), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x82y67     80'h00_0060_00_0000_0C08_FFB3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a600_4 ( .OUT(na600_2), .IN1(1'b0), .IN2(~na1952_2), .IN3(na1329_1), .IN4(~na11_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x83y60     80'h00_0018_00_0000_0C88_BAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a603_1 ( .OUT(na603_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b0), .IN7(na521_1), .IN8(~na604_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x88y50     80'h00_0018_00_0040_0A33_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a604_1 ( .OUT(na604_1), .IN1(na1064_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1555_2), .IN6(~na1149_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y74     80'h00_0018_00_0000_0888_F5DC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a608_1 ( .OUT(na608_1), .IN1(1'b0), .IN2(na101_1), .IN3(~na331_1), .IN4(na11_1), .IN5(~na1547_1), .IN6(1'b0), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x98y47     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a611_1 ( .OUT(na611_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b0), .IN7(na612_1), .IN8(na1563_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y47     80'h00_0018_00_0000_0C88_15FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a612_1 ( .OUT(na612_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na613_1), .IN6(1'b1), .IN7(~na2031_2), .IN8(~na1065_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x87y47     80'h00_0018_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a613_1 ( .OUT(na613_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na510_1), .IN4(1'b1), .IN5(1'b0), .IN6(na509_1), .IN7(1'b0), .IN8(na511_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x87y60     80'h00_0018_00_0000_0EEE_CDCE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a616_1 ( .OUT(na616_1), .IN1(na1577_1), .IN2(na625_1), .IN3(1'b0), .IN4(na2115_2), .IN5(~na1581_1), .IN6(na1568_1), .IN7(1'b0),
                     .IN8(na1582_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x84y68     80'h00_0078_00_0000_0C88_C58F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a617_1 ( .OUT(na617_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na587_1), .IN6(1'b1), .IN7(1'b1), .IN8(na102_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a617_4 ( .OUT(na617_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1576_1), .IN4(na102_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x72y51     80'h00_0018_00_0040_0A76_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a620_1 ( .OUT(na620_1), .IN1(1'b1), .IN2(~na2087_2), .IN3(1'b1), .IN4(na24_1), .IN5(na85_1), .IN6(~na2074_2), .IN7(~na1337_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x91y52     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a625_1 ( .OUT(na625_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b0), .IN7(na612_1), .IN8(na1580_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x83y68     80'h00_0018_00_0000_0C88_54FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a628_1 ( .OUT(na628_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1515_1), .IN6(na101_1), .IN7(~na572_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x95y51     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a632_1 ( .OUT(na632_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b0), .IN7(na612_1), .IN8(na1588_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x85y73     80'h00_0018_00_0000_0C88_43FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a635_1 ( .OUT(na635_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na560_1), .IN7(~na1501_1), .IN8(na1907_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x94y52     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a639_1 ( .OUT(na639_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b0), .IN7(na612_1), .IN8(na1596_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x88y53     80'h00_0018_00_0000_0EEE_AAEB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a641_1 ( .OUT(na641_1), .IN1(na830_1), .IN2(~na1607_1), .IN3(na1599_2), .IN4(na646_1), .IN5(na1608_1), .IN6(1'b0), .IN7(na1599_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x83y64     80'h00_0018_00_0000_0C88_43FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a642_1 ( .OUT(na642_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na548_1), .IN7(~na1489_1), .IN8(na1907_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x91y63     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a643_1 ( .OUT(na643_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1494_1), .IN6(na1952_2), .IN7(1'b0), .IN8(na102_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x92y50     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a646_1 ( .OUT(na646_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b0), .IN7(na612_1), .IN8(na1606_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x83y73     80'h00_0018_00_0000_0888_DF7C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a648_1 ( .OUT(na648_1), .IN1(1'b0), .IN2(na101_1), .IN3(~na1479_1), .IN4(~na11_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na536_1),
                     .IN8(na11_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x94y67     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a649_1 ( .OUT(na649_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1481_1), .IN6(na1952_2), .IN7(1'b0), .IN8(na102_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x82y71     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a652_1 ( .OUT(na652_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b0), .IN7(na612_1), .IN8(na1614_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x88y56     80'h00_0018_00_0000_0EEE_AAEE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a655_1 ( .OUT(na655_1), .IN1(na662_2), .IN2(na1624_1), .IN3(na1619_1), .IN4(na660_1), .IN5(na662_1), .IN6(1'b0), .IN7(na1619_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x82y59     80'h00_0018_00_0000_0888_7B7D
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a656_1 ( .OUT(na656_1), .IN1(~na1910_2), .IN2(na1470_1), .IN3(~na1623_1), .IN4(~na102_1), .IN5(na1961_2), .IN6(~na101_1),
                     .IN7(~na834_1), .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x92y52     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a660_1 ( .OUT(na660_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b0), .IN7(na612_1), .IN8(na1626_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x89y67     80'h00_0078_00_0000_0C88_ACCA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a662_1 ( .OUT(na662_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na942_1), .IN7(na346_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a662_4 ( .OUT(na662_2), .IN1(na917_2), .IN2(1'b1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x87y74     80'h00_0018_00_0000_0888_DF7C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a664_1 ( .OUT(na664_1), .IN1(1'b0), .IN2(na101_1), .IN3(~na1460_1), .IN4(~na11_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na495_1),
                     .IN8(na11_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x96y69     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a665_1 ( .OUT(na665_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1630_2), .IN6(na1952_2), .IN7(1'b0), .IN8(na102_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x95y50     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a669_1 ( .OUT(na669_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b0), .IN7(na612_1), .IN8(na1635_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x84y54     80'h00_0018_00_0000_0888_77BD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a671_1 ( .OUT(na671_1), .IN1(~na1341_2), .IN2(na1643_2), .IN3(na672_1), .IN4(~na350_1), .IN5(~na1062_2), .IN6(~na567_1),
                     .IN7(~na1045_2), .IN8(~na350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x90y63     80'h00_0018_00_0000_0888_7B7B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a672_1 ( .OUT(na672_1), .IN1(na1440_1), .IN2(~na1911_2), .IN3(~na1642_1), .IN4(~na102_1), .IN5(na496_1), .IN6(~na101_1),
                     .IN7(~na839_1), .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y54     80'h00_0018_00_0000_0888_77BD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a677_1 ( .OUT(na677_1), .IN1(~na1341_2), .IN2(na1652_1), .IN3(na678_1), .IN4(~na350_1), .IN5(~na1077_2), .IN6(~na567_1),
                     .IN7(~na868_1), .IN8(~na350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x80y63     80'h00_0018_00_0000_0888_777B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a678_1 ( .OUT(na678_1), .IN1(na1431_1), .IN2(~na1911_2), .IN3(~na1651_1), .IN4(~na102_1), .IN5(~na1957_2), .IN6(~na101_1),
                     .IN7(~na841_1), .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x83y54     80'h00_0018_00_0000_0888_77BD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a683_1 ( .OUT(na683_1), .IN1(~na1341_2), .IN2(na1662_1), .IN3(na1657_1), .IN4(~na350_1), .IN5(~na1077_1), .IN6(~na567_1),
                     .IN7(~na1047_2), .IN8(~na350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x84y65     80'h00_0078_00_0000_0C88_AC3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a684_1 ( .OUT(na684_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na101_1), .IN7(na460_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a684_4 ( .OUT(na684_2), .IN1(1'b1), .IN2(na1909_2), .IN3(1'b1), .IN4(~na688_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x72y50     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a687_1 ( .OUT(na687_1), .IN1(~na2111_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1894_2), .IN5(na85_1), .IN6(~na2074_2), .IN7(~na1337_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x68y76     80'h00_0018_00_0040_0C55_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a688_1 ( .OUT(na688_1), .IN1(~na970_1), .IN2(1'b0), .IN3(~na1002_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na335_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x71y63     80'h00_0018_00_0000_0C88_C2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a689_1 ( .OUT(na689_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na84_1), .IN6(~na33_1), .IN7(1'b1), .IN8(na1514_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y56     80'h00_0018_00_0000_0888_77BD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a693_1 ( .OUT(na693_1), .IN1(~na1341_2), .IN2(na1676_2), .IN3(na1667_1), .IN4(~na350_1), .IN5(~na1079_2), .IN6(~na567_1),
                     .IN7(~na1968_2), .IN8(~na350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x74y47     80'h00_0018_00_0040_0A76_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a695_1 ( .OUT(na695_1), .IN1(na34_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1510_2), .IN5(na85_1), .IN6(~na2074_2), .IN7(~na1337_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x83y62     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a698_1 ( .OUT(na698_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2081_2), .IN6(na1952_2), .IN7(1'b0), .IN8(na102_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x83y55     80'h00_0018_00_0000_0888_7D77
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a702_1 ( .OUT(na702_1), .IN1(~na1079_1), .IN2(~na567_1), .IN3(~na1681_1), .IN4(~na350_1), .IN5(~na1341_2), .IN6(na1687_2),
                     .IN7(~na1049_2), .IN8(~na350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x72y49     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a706_1 ( .OUT(na706_1), .IN1(~na2110_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1895_2), .IN5(na85_1), .IN6(~na2074_2), .IN7(~na1337_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x80y77     80'h00_0018_00_0040_0CAA_CF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a707_1 ( .OUT(na707_1), .IN1(1'b0), .IN2(~na972_1), .IN3(1'b0), .IN4(~na1004_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na335_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x76y62     80'h00_0018_00_0000_0C88_A4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a708_1 ( .OUT(na708_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na35_1), .IN6(na1906_2), .IN7(na1509_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x77y65     80'h00_0018_00_0000_0888_77BD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a711_1 ( .OUT(na711_1), .IN1(~na1341_2), .IN2(na1698_1), .IN3(na1692_1), .IN4(~na350_1), .IN5(~na1081_2), .IN6(~na567_1),
                     .IN7(~na872_1), .IN8(~na350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x88y65     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a714_1 ( .OUT(na714_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2079_2), .IN6(na1952_2), .IN7(1'b0), .IN8(na102_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y56     80'h00_0018_00_0000_0888_7DB5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a718_1 ( .OUT(na718_1), .IN1(~na726_1), .IN2(1'b0), .IN3(na719_1), .IN4(~na350_1), .IN5(~na1341_2), .IN6(na1712_1), .IN7(~na1051_1),
                     .IN8(~na350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x84y57     80'h00_0018_00_0000_0888_4F1C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a719_1 ( .OUT(na719_1), .IN1(1'b1), .IN2(na1708_1), .IN3(~na1705_1), .IN4(~na721_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1705_2),
                     .IN8(na1703_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x72y52     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a721_1 ( .OUT(na721_1), .IN1(~na2108_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1897_2), .IN5(na85_1), .IN6(~na2074_2), .IN7(~na1337_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x79y57     80'h00_0018_00_0000_0C88_48FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a726_1 ( .OUT(na726_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1053_2), .IN6(na1940_2), .IN7(~na1055_2),
                     .IN8(na5_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y57     80'h00_0018_00_0000_0888_77BD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a727_1 ( .OUT(na727_1), .IN1(~na1341_2), .IN2(na1721_2), .IN3(na1715_1), .IN4(~na350_1), .IN5(~na1964_2), .IN6(~na1063_2),
                     .IN7(~na1969_2), .IN8(~na350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x84y75     80'h00_0018_00_0000_0C88_ECFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a728_1 ( .OUT(na728_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na101_1), .IN7(na1967_2), .IN8(na298_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y56     80'h00_0018_00_0040_0A7F_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a731_1 ( .OUT(na731_1), .IN1(na38_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1497_2), .IN5(~na84_1), .IN6(~na1904_2), .IN7(~na83_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x71y63     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a732_4 ( .OUT(na732_2), .IN1(na1720_1), .IN2(1'b1), .IN3(1'b1), .IN4(na102_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x87y54     80'h00_0018_00_0000_0888_3FD3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a736_1 ( .OUT(na736_1), .IN1(1'b0), .IN2(~na1228_2), .IN3(~na240_2), .IN4(na1056_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x61y65     80'h00_0018_00_0000_0888_FB5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a737_1 ( .OUT(na737_1), .IN1(1'b0), .IN2(na738_1), .IN3(~na510_2), .IN4(1'b0), .IN5(na1064_1), .IN6(~na1982_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x67y50     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a738_1 ( .OUT(na738_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2021_2), .IN7(na240_2), .IN8(na44_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x61y67     80'h00_0018_00_0000_0888_FB5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a739_1 ( .OUT(na739_1), .IN1(1'b0), .IN2(na738_1), .IN3(~na510_1), .IN4(1'b0), .IN5(na1064_1), .IN6(~na1982_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x61y68     80'h00_0018_00_0000_0888_FE5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a740_1 ( .OUT(na740_1), .IN1(1'b0), .IN2(na738_1), .IN3(~na510_2), .IN4(1'b0), .IN5(na1064_1), .IN6(na1982_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x61y71     80'h00_0018_00_0000_0888_FE5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a741_1 ( .OUT(na741_1), .IN1(1'b0), .IN2(na738_1), .IN3(~na510_1), .IN4(1'b0), .IN5(na1064_1), .IN6(na1982_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x73y69     80'h00_0018_00_0040_0C85_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a774_1 ( .OUT(na774_1), .IN1(na274_1), .IN2(1'b0), .IN3(na272_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na4_1), .IN7(1'b1), .IN8(na7_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y59     80'h00_0018_00_0040_0A3B_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a775_1 ( .OUT(na775_1), .IN1(~na774_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1868_2), .IN5(~na273_1), .IN6(~na275_1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x80y72     80'h00_0018_00_0040_0C23_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a776_1 ( .OUT(na776_1), .IN1(na775_1), .IN2(~na276_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na8_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x85y75     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a777_1 ( .OUT(na777_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1730_1), .IN7(1'b1), .IN8(na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x73y56     80'h00_0018_00_0040_0C8A_3F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a778_1 ( .OUT(na778_1), .IN1(1'b0), .IN2(na1731_1), .IN3(1'b0), .IN4(~na1243_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1065_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x78y74     80'h00_0018_00_0040_0C53_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a780_1 ( .OUT(na780_1), .IN1(~na355_1), .IN2(na353_1), .IN3(1'b1), .IN4(1'b0), .IN5(1'b1), .IN6(~na8_1), .IN7(1'b1), .IN8(~na7_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x78y72     80'h00_0018_00_0040_0AA1_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a781_1 ( .OUT(na781_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b1), .IN4(~na780_1), .IN5(1'b1), .IN6(na356_1), .IN7(1'b0), .IN8(na354_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y81     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a782_1 ( .OUT(na782_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1735_2), .IN6(na357_1), .IN7(1'b0), .IN8(na11_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y55     80'h00_0018_00_0040_0A76_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a783_1 ( .OUT(na783_1), .IN1(1'b1), .IN2(~na2104_2), .IN3(1'b1), .IN4(na7_1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y61     80'h00_0018_00_0040_0A76_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a785_1 ( .OUT(na785_1), .IN1(1'b1), .IN2(~na2102_2), .IN3(1'b1), .IN4(na1873_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x72y57     80'h00_0018_00_0000_0EEE_ADC5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a787_1 ( .OUT(na787_1), .IN1(~na1376_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1379_2), .IN5(~na1376_2), .IN6(na1738_2), .IN7(na1375_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y57     80'h00_0018_00_0040_0A76_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a788_1 ( .OUT(na788_1), .IN1(1'b1), .IN2(~na2101_2), .IN3(na10_1), .IN4(1'b1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x67y59     80'h00_0018_00_0040_0A76_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a789_1 ( .OUT(na789_1), .IN1(1'b1), .IN2(~na2098_2), .IN3(1'b1), .IN4(na1878_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y49     80'h00_0018_00_0040_0A76_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a790_1 ( .OUT(na790_1), .IN1(1'b1), .IN2(~na2097_2), .IN3(1'b1), .IN4(na1879_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x82y53     80'h00_0018_00_0000_0EEE_5AAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a792_1 ( .OUT(na792_1), .IN1(na1439_2), .IN2(na1435_1), .IN3(na493_1), .IN4(1'b0), .IN5(na1741_2), .IN6(1'b0), .IN7(~na1438_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x78y48     80'h00_0018_00_0040_0A76_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a793_1 ( .OUT(na793_1), .IN1(1'b1), .IN2(~na2096_2), .IN3(na1880_2), .IN4(1'b1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x82y55     80'h00_0018_00_0000_0EEE_A3CB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a794_1 ( .OUT(na794_1), .IN1(na1453_2), .IN2(~na1450_1), .IN3(1'b0), .IN4(na1449_1), .IN5(1'b0), .IN6(~na1450_2), .IN7(na1743_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x90y56     80'h00_0018_00_0000_0888_BF73
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a795_1 ( .OUT(na795_1), .IN1(1'b0), .IN2(~na494_2), .IN3(~na1448_1), .IN4(~na102_1), .IN5(1'b1), .IN6(1'b1), .IN7(na1958_2),
                     .IN8(~na102_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x68y60     80'h00_0018_00_0040_0C15_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a796_1 ( .OUT(na796_1), .IN1(~na1745_1), .IN2(1'b0), .IN3(na794_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na795_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x76y51     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a797_1 ( .OUT(na797_1), .IN1(~na2095_2), .IN2(1'b1), .IN3(1'b1), .IN4(na15_1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x77y51     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a800_1 ( .OUT(na800_1), .IN1(~na2094_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1882_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x84y55     80'h00_0018_00_0000_0EEE_D0CE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a802_1 ( .OUT(na802_1), .IN1(na1477_1), .IN2(na533_2), .IN3(1'b0), .IN4(na1473_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na1476_1),
                     .IN8(na1750_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y54     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a803_1 ( .OUT(na803_1), .IN1(~na2093_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1883_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x85y54     80'h00_0018_00_0000_0EEE_5AAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a805_1 ( .OUT(na805_1), .IN1(na1753_2), .IN2(na1485_1), .IN3(na1487_2), .IN4(1'b0), .IN5(na1483_1), .IN6(1'b0), .IN7(~na1486_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y53     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a806_1 ( .OUT(na806_1), .IN1(~na2092_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1884_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x85y55     80'h00_0018_00_0000_0EEE_AD0E
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a809_1 ( .OUT(na809_1), .IN1(na1757_1), .IN2(na1756_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1499_1), .IN6(na1500_2), .IN7(na1498_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x70y49     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a810_1 ( .OUT(na810_1), .IN1(~na2091_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1885_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x87y58     80'h00_0018_00_0000_0EEE_E5AB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a812_1 ( .OUT(na812_1), .IN1(na1512_2), .IN2(~na1507_1), .IN3(na1760_1), .IN4(1'b0), .IN5(~na1511_1), .IN6(1'b0), .IN7(na1506_2),
                     .IN8(na1508_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x78y53     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a813_1 ( .OUT(na813_1), .IN1(~na2090_2), .IN2(1'b1), .IN3(1'b1), .IN4(na20_1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x72y63     80'h00_0018_00_0040_0A76_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a815_1 ( .OUT(na815_1), .IN1(na21_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1452_1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x78y55     80'h00_0018_00_0040_0A76_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a817_1 ( .OUT(na817_1), .IN1(na22_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1447_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x75y55     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a819_1 ( .OUT(na819_1), .IN1(~na2089_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1887_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x87y59     80'h00_0018_00_0000_0EEE_E3E5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a821_1 ( .OUT(na821_1), .IN1(~na1564_1), .IN2(1'b0), .IN3(na1565_2), .IN4(na1766_2), .IN5(1'b0), .IN6(~na1566_1), .IN7(na611_1),
                     .IN8(na1567_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x71y53     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a822_1 ( .OUT(na822_1), .IN1(~na2086_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1889_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x88y62     80'h00_0018_00_0000_0EEE_DEE0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a824_1 ( .OUT(na824_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1585_2), .IN4(na1769_2), .IN5(na632_1), .IN6(na1590_2), .IN7(~na1589_1),
                     .IN8(na1769_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x72y55     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a825_1 ( .OUT(na825_1), .IN1(~na2085_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1890_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x87y61     80'h00_0018_00_0000_0EEE_EB0E
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a827_1 ( .OUT(na827_1), .IN1(na1772_1), .IN2(na1593_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1772_2), .IN6(~na1597_1), .IN7(na1598_2),
                     .IN8(na639_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y49     80'h00_0018_00_0040_0A76_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a828_1 ( .OUT(na828_1), .IN1(na27_1), .IN2(1'b1), .IN3(~na1525_1), .IN4(1'b1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y55     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a830_1 ( .OUT(na830_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1775_1), .IN7(1'b1), .IN8(na350_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y49     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a831_1 ( .OUT(na831_1), .IN1(~na2114_2), .IN2(1'b1), .IN3(1'b1), .IN4(na28_1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x87y53     80'h00_0018_00_0000_0EEE_BACB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a833_1 ( .OUT(na833_1), .IN1(na1616_1), .IN2(~na1615_2), .IN3(1'b0), .IN4(na1778_2), .IN5(na1618_1), .IN6(1'b0), .IN7(na652_1),
                     .IN8(~na1617_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y51     80'h00_0018_00_0040_0A76_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a834_1 ( .OUT(na834_1), .IN1(na29_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1519_1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x81y51     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a836_1 ( .OUT(na836_1), .IN1(~na2113_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1892_2), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x88y59     80'h00_0018_00_0000_0EEE_BCEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a838_1 ( .OUT(na838_1), .IN1(1'b0), .IN2(na2116_2), .IN3(na1782_2), .IN4(na1632_2), .IN5(1'b0), .IN6(na669_1), .IN7(na1637_1),
                     .IN8(~na1636_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x78y49     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a839_1 ( .OUT(na839_1), .IN1(~na2112_2), .IN2(1'b1), .IN3(1'b1), .IN4(na31_1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y53     80'h00_0018_00_0040_0A76_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a841_1 ( .OUT(na841_1), .IN1(na32_1), .IN2(1'b1), .IN3(~na1516_2), .IN4(1'b1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x86y63     80'h00_0018_00_0040_0A76_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a843_1 ( .OUT(na843_1), .IN1(~na2109_2), .IN2(1'b1), .IN3(1'b1), .IN4(na36_1), .IN5(na1064_1), .IN6(~na1063_1), .IN7(~na2029_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x87y62     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a845_1 ( .OUT(na845_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na788_1), .IN6(na1788_2), .IN7(1'b0), .IN8(na1065_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x86y51     80'h00_0018_00_0000_0EEE_AAE3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a847_1 ( .OUT(na847_1), .IN1(1'b0), .IN2(~na1394_2), .IN3(na1790_2), .IN4(na1390_1), .IN5(na1391_2), .IN6(1'b0), .IN7(na1395_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x89y59     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a848_1 ( .OUT(na848_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na789_1), .IN6(na1793_1), .IN7(1'b0), .IN8(na1065_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x83y51     80'h00_0018_00_0000_0EEE_0BAB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a850_1 ( .OUT(na850_1), .IN1(na1426_2), .IN2(~na1421_2), .IN3(na1795_1), .IN4(1'b0), .IN5(na1422_2), .IN6(~na1421_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y56     80'h00_FE60_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a853_1 ( .OUT(na853_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na853_1),
                     .CINX(1'b0), .CINY1(na882_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a853_2 ( .OUT(na853_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na853_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a853_4 ( .OUT(na853_2), .COUTY1(na853_4), .IN1(na1033_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na853_1), .CINX(1'b0), .CINY1(na882_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y57     80'h00_FE60_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a855_1 ( .OUT(na855_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na855_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na853_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a855_2 ( .OUT(na855_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na855_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a855_4 ( .OUT(na855_2), .COUTY1(na855_4), .IN1(1'b1), .IN2(na1035_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na855_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na853_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y58     80'h00_FE60_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a857_1 ( .OUT(na857_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na857_1),
                     .CINX(1'b0), .CINY1(na855_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a857_2 ( .OUT(na857_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na857_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a857_4 ( .OUT(na857_2), .COUTY1(na857_4), .IN1(na1037_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na857_1), .CINX(1'b0), .CINY1(na855_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y59     80'h00_FE60_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a859_1 ( .OUT(na859_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na859_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na857_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a859_2 ( .OUT(na859_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na859_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a859_4 ( .OUT(na859_2), .COUTY1(na859_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1039_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na859_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na857_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y60     80'h00_FE60_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a861_1 ( .OUT(na861_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na861_1),
                     .CINX(1'b0), .CINY1(na859_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a861_2 ( .OUT(na861_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na861_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a861_4 ( .OUT(na861_2), .COUTY1(na861_4), .IN1(na1041_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na861_1), .CINX(1'b0), .CINY1(na859_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y51     80'h00_FE60_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a862_1 ( .OUT(na862_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1023_2), .IN7(na862_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na907_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a862_2 ( .OUT(na862_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na862_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a862_4 ( .OUT(na862_2), .COUTY1(na862_4), .IN1(1'b1), .IN2(na1023_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1023_2),
                     .IN7(na862_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na907_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y61     80'h00_FE60_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a864_1 ( .OUT(na864_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na864_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na861_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a864_2 ( .OUT(na864_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na864_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a864_4 ( .OUT(na864_2), .COUTY1(na864_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1043_1), .IN5(1'b0), .IN6(1'b0), .IN7(na864_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na861_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y62     80'h00_FE60_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a866_1 ( .OUT(na866_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na866_1),
                     .CINX(1'b0), .CINY1(na864_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a866_2 ( .OUT(na866_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na866_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a866_4 ( .OUT(na866_2), .COUTY1(na866_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1045_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na866_1), .CINX(1'b0), .CINY1(na864_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y63     80'h00_FE60_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a868_1 ( .OUT(na868_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na868_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na866_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a868_2 ( .OUT(na868_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na868_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a868_4 ( .OUT(na868_2), .COUTY1(na868_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1047_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na868_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na866_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y64     80'h00_FE60_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a870_1 ( .OUT(na870_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na870_1),
                     .CINX(1'b0), .CINY1(na868_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a870_2 ( .OUT(na870_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na870_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a870_4 ( .OUT(na870_2), .COUTY1(na870_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1049_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na870_1), .CINX(1'b0), .CINY1(na868_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y65     80'h00_FE60_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a872_1 ( .OUT(na872_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na872_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na870_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a872_2 ( .OUT(na872_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na872_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a872_4 ( .OUT(na872_2), .COUTY1(na872_4), .IN1(1'b0), .IN2(1'b0), .IN3(na1051_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na872_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na870_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF/D///      x96y66     80'h00_FE00_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a875_1 ( .OUT(na875_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na875_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na872_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a875_2 ( .OUT(na875_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na875_1_i) );
// C_ADDF2/D//ADDF2/      x96y52     80'h00_FE60_00_0020_0C66_C00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a876_1 ( .OUT(na876_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na876_1),
                     .CINX(1'b0), .CINY1(na862_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a876_2 ( .OUT(na876_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na876_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a876_4 ( .OUT(na876_2), .COUTY1(na876_4), .IN1(1'b1), .IN2(na1025_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na876_1), .CINX(1'b0), .CINY1(na862_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y53     80'h00_FE60_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a878_1 ( .OUT(na878_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na878_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na876_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a878_2 ( .OUT(na878_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na878_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a878_4 ( .OUT(na878_2), .COUTY1(na878_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1027_2), .IN5(1'b0), .IN6(1'b0), .IN7(na878_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na876_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y54     80'h00_FE60_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a880_1 ( .OUT(na880_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na880_1),
                     .CINX(1'b0), .CINY1(na878_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a880_2 ( .OUT(na880_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na880_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a880_4 ( .OUT(na880_2), .COUTY1(na880_4), .IN1(na1029_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na880_1), .CINX(1'b0), .CINY1(na878_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x96y55     80'h00_FE60_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a882_1 ( .OUT(na882_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na882_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na880_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a882_2 ( .OUT(na882_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na882_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a882_4 ( .OUT(na882_2), .COUTY1(na882_4), .IN1(na1031_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na882_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na880_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x78y57     80'h00_0018_00_0010_0666_20A8
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a883_1 ( .OUT(na883_1), .COUTY1(na883_4), .IN1(na1058_1), .IN2(na2021_2), .IN3(na1496_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0),
                     .IN7(na2023_2), .IN8(~na1056_1), .CINX(1'b0), .CINY1(na1009_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x78y65     80'h00_0078_00_0020_0C66_CCAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a885_1 ( .OUT(na885_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1063_2), .IN7(1'b1), .IN8(na1459_2),
                     .CINX(1'b0), .CINY1(na906_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a885_4 ( .OUT(na885_2), .COUTY1(na885_4), .IN1(1'b1), .IN2(na1063_2), .IN3(na1455_1), .IN4(1'b1), .IN5(1'b1), .IN6(na1063_2),
                     .IN7(1'b1), .IN8(na1459_2), .CINX(1'b0), .CINY1(na906_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x78y66     80'h00_0078_00_0020_0C66_ACCC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a887_1 ( .OUT(na887_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1063_2), .IN7(na1454_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na885_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a887_4 ( .OUT(na887_2), .COUTY1(na887_4), .IN1(1'b1), .IN2(na1063_2), .IN3(1'b1), .IN4(na1452_1), .IN5(1'b1), .IN6(na1063_2),
                     .IN7(na1454_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na885_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x78y67     80'h00_0078_00_0020_0C66_CCAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a889_1 ( .OUT(na889_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1063_2), .IN7(1'b1), .IN8(na1447_2),
                     .CINX(1'b0), .CINY1(na887_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a889_4 ( .OUT(na889_2), .COUTY1(na889_4), .IN1(1'b1), .IN2(na1063_2), .IN3(na1442_1), .IN4(1'b1), .IN5(1'b1), .IN6(na1063_2),
                     .IN7(1'b1), .IN8(na1447_2), .CINX(1'b0), .CINY1(na887_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x78y68     80'h00_0078_00_0020_0C66_ACCC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a891_1 ( .OUT(na891_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1063_2), .IN7(na1436_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na889_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a891_4 ( .OUT(na891_2), .COUTY1(na891_4), .IN1(1'b1), .IN2(na1063_2), .IN3(1'b1), .IN4(na1433_1), .IN5(1'b1), .IN6(na1063_2),
                     .IN7(na1436_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na889_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x78y69     80'h00_0078_00_0020_0C66_CCAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a893_1 ( .OUT(na893_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1063_2), .IN7(1'b1), .IN8(na1430_2),
                     .CINX(1'b0), .CINY1(na891_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a893_4 ( .OUT(na893_2), .COUTY1(na893_4), .IN1(1'b1), .IN2(na1063_2), .IN3(na1525_1), .IN4(1'b1), .IN5(1'b1), .IN6(na1063_2),
                     .IN7(1'b1), .IN8(na1430_2), .CINX(1'b0), .CINY1(na891_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x78y58     80'h00_0018_00_0010_0666_20A8
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a894_1 ( .OUT(na894_1), .COUTY1(na894_4), .IN1(na1059_1), .IN2(na2021_2), .IN3(na1493_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0),
                     .IN7(na2024_2), .IN8(~na1056_1), .CINX(1'b0), .CINY1(na883_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x78y70     80'h00_0078_00_0020_0C66_ACCC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a896_1 ( .OUT(na896_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1063_2), .IN7(na1520_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na893_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a896_4 ( .OUT(na896_2), .COUTY1(na896_4), .IN1(1'b1), .IN2(na1063_2), .IN3(1'b1), .IN4(na1519_1), .IN5(1'b1), .IN6(na1063_2),
                     .IN7(na1520_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na893_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x78y71     80'h00_0018_00_0010_0666_00CC
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a898_1 ( .OUT(na898_1), .IN1(1'b1), .IN2(na1063_2), .IN3(1'b1), .IN4(na1518_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na896_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x78y59     80'h00_0018_00_0010_0666_208C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a899_1 ( .OUT(na899_1), .COUTY1(na899_4), .IN1(1'b1), .IN2(na2102_2), .IN3(na1060_1), .IN4(na1056_1), .IN5(1'b0), .IN6(1'b0),
                     .IN7(na1060_2), .IN8(~na1056_1), .CINX(1'b0), .CINY1(na894_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x78y60     80'h00_0018_00_0010_0666_20C8
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a900_1 ( .OUT(na900_1), .COUTY1(na900_4), .IN1(na1061_1), .IN2(na2021_2), .IN3(1'b1), .IN4(na1491_2), .IN5(1'b0), .IN6(1'b0),
                     .IN7(na2027_2), .IN8(~na1056_1), .CINX(1'b0), .CINY1(na899_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x78y61     80'h00_0018_00_0010_0666_20A8
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a901_1 ( .OUT(na901_1), .COUTY1(na901_4), .IN1(na1062_1), .IN2(na2021_2), .IN3(na1484_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0),
                     .IN7(na2028_2), .IN8(~na1056_1), .CINX(1'b0), .CINY1(na900_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x78y62     80'h00_0078_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a902_1 ( .OUT(na902_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1077_2), .IN6(1'b1), .IN7(na1480_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na901_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a902_4 ( .OUT(na902_2), .COUTY1(na902_4), .IN1(na1077_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1478_1), .IN5(na1077_2), .IN6(1'b1),
                     .IN7(na1480_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na901_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x78y63     80'h00_0078_00_0020_0C66_CAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a904_1 ( .OUT(na904_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1079_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1475_2),
                     .CINX(1'b0), .CINY1(na902_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a904_4 ( .OUT(na904_2), .COUTY1(na904_4), .IN1(na1079_1), .IN2(1'b1), .IN3(na1474_1), .IN4(1'b1), .IN5(na1079_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na1475_2), .CINX(1'b0), .CINY1(na902_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x78y64     80'h00_0078_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a906_1 ( .OUT(na906_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1081_2), .IN6(1'b1), .IN7(na1468_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na904_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a906_4 ( .OUT(na906_2), .COUTY1(na906_4), .IN1(na1081_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1463_1), .IN5(na1081_2), .IN6(1'b1),
                     .IN7(na1468_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na904_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x96y50     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a907_2 ( .OUT(na907_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a907_6 ( .COUTY1(na907_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na907_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x95y67     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a909_1 ( .OUT(na909_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na260_2),
                     .CINX(1'b0), .CINY1(na928_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a909_4 ( .OUT(na909_2), .COUTY1(na909_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na260_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na260_2), .CINX(1'b0), .CINY1(na928_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x95y68     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a911_1 ( .OUT(na911_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na262_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na909_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a911_4 ( .OUT(na911_2), .COUTY1(na911_4), .IN1(1'b1), .IN2(na262_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na262_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na909_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x95y69     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a913_1 ( .OUT(na913_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na264_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na911_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a913_4 ( .OUT(na913_2), .COUTY1(na913_4), .IN1(1'b1), .IN2(na264_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na264_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na911_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x95y70     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a915_1 ( .OUT(na915_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na266_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na913_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a915_4 ( .OUT(na915_2), .COUTY1(na915_4), .IN1(1'b1), .IN2(na266_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na266_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na913_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x95y71     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a917_1 ( .OUT(na917_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na268_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na915_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a917_4 ( .OUT(na917_2), .COUTY1(na917_4), .IN1(1'b1), .IN2(na268_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na268_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na915_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x95y62     80'h00_0078_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a918_1 ( .OUT(na918_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na249_1), .IN7(1'b1), .IN8(na250_2),
                     .CINX(1'b0), .CINY1(na1222_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a918_4 ( .OUT(na918_2), .COUTY1(na918_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na250_1), .IN5(1'b1), .IN6(na249_1), .IN7(1'b1),
                     .IN8(na250_2), .CINX(1'b0), .CINY1(na1222_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x95y72     80'h00_0018_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a920_1 ( .OUT(na920_1), .IN1(1'b1), .IN2(na269_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na917_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x95y63     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a922_1 ( .OUT(na922_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na252_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na918_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a922_4 ( .OUT(na922_2), .COUTY1(na922_4), .IN1(1'b1), .IN2(na252_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na252_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na918_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x95y64     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a924_1 ( .OUT(na924_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na254_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na922_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a924_4 ( .OUT(na924_2), .COUTY1(na924_4), .IN1(1'b1), .IN2(na254_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na254_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na922_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x95y65     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a926_1 ( .OUT(na926_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na256_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na924_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a926_4 ( .OUT(na926_2), .COUTY1(na926_4), .IN1(1'b1), .IN2(na256_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na256_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na924_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x95y66     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a928_1 ( .OUT(na928_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na258_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na926_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a928_4 ( .OUT(na928_2), .COUTY1(na928_4), .IN1(1'b1), .IN2(na258_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na258_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na926_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y56     80'h00_0018_00_0010_0666_08A2
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a929_1 ( .OUT(na929_1), .COUTY1(na929_4), .IN1(na1223_2), .IN2(~na1054_1), .IN3(na247_2), .IN4(1'b1), .IN5(na1059_2), .IN6(na1054_1),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1232_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y63     80'h00_0018_00_0010_0666_08C2
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a930_1 ( .OUT(na930_1), .COUTY1(na930_4), .IN1(na1227_2), .IN2(~na1054_1), .IN3(1'b1), .IN4(na1918_2), .IN5(na1058_2), .IN6(na1054_1),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na950_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y64     80'h00_0018_00_0010_0666_08C4
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a931_1 ( .OUT(na931_1), .COUTY1(na931_4), .IN1(~na45_1), .IN2(na1063_1), .IN3(1'b1), .IN4(na1917_2), .IN5(na45_1), .IN6(na1063_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na930_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y65     80'h00_0018_00_0010_0666_08C2
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a932_1 ( .OUT(na932_1), .COUTY1(na932_4), .IN1(na1064_1), .IN2(~na1900_2), .IN3(1'b1), .IN4(na260_2), .IN5(na45_1), .IN6(na1063_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na931_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y66     80'h00_0018_00_0010_0666_084C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a933_1 ( .OUT(na933_1), .COUTY1(na933_4), .IN1(1'b1), .IN2(na1919_2), .IN3(~na1901_2), .IN4(na1065_2), .IN5(na45_1), .IN6(na1063_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na932_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y67     80'h00_0018_00_0010_0666_08C4
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a934_1 ( .OUT(na934_1), .COUTY1(na934_4), .IN1(~na45_1), .IN2(na2034_2), .IN3(1'b1), .IN4(na1922_2), .IN5(na45_1), .IN6(na1063_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na933_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y68     80'h00_0018_00_0010_0666_08C4
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a935_1 ( .OUT(na935_1), .COUTY1(na935_4), .IN1(~na45_1), .IN2(na2035_2), .IN3(1'b1), .IN4(na1921_2), .IN5(na45_1), .IN6(na1063_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na934_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y69     80'h00_0018_00_0010_0666_08C4
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a936_1 ( .OUT(na936_1), .COUTY1(na936_4), .IN1(~na45_1), .IN2(na2036_2), .IN3(1'b1), .IN4(na1924_2), .IN5(na45_1), .IN6(na1063_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na935_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y70     80'h00_0018_00_0010_0666_08C4
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a937_1 ( .OUT(na937_1), .COUTY1(na937_4), .IN1(~na45_1), .IN2(na2037_2), .IN3(1'b1), .IN4(na1923_2), .IN5(na45_1), .IN6(na1063_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na936_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y71     80'h00_0018_00_0010_0666_08C4
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a938_1 ( .OUT(na938_1), .COUTY1(na938_4), .IN1(~na45_1), .IN2(na2038_2), .IN3(1'b1), .IN4(na1926_2), .IN5(na45_1), .IN6(na1063_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na937_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y72     80'h00_0018_00_0010_0666_80C4
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a939_1 ( .OUT(na939_1), .COUTY1(na939_4), .IN1(~na1869_2), .IN2(na1063_2), .IN3(1'b1), .IN4(na1925_2), .IN5(1'b0), .IN6(1'b0),
                     .IN7(na2023_2), .IN8(na5_2), .CINX(1'b0), .CINY1(na938_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y57     80'h00_0018_00_0010_0666_08C2
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a940_1 ( .OUT(na940_1), .COUTY1(na940_4), .IN1(na1224_1), .IN2(~na1054_1), .IN3(1'b1), .IN4(na250_2), .IN5(na2025_2), .IN6(na1054_1),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na929_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y73     80'h00_0018_00_0010_0666_80C4
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a941_1 ( .OUT(na941_1), .COUTY1(na941_4), .IN1(~na1869_2), .IN2(na1063_2), .IN3(1'b1), .IN4(na1928_2), .IN5(1'b0), .IN6(1'b0),
                     .IN7(na2024_2), .IN8(na5_2), .CINX(1'b0), .CINY1(na939_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y74     80'h00_0018_00_0010_0666_80C4
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a942_1 ( .OUT(na942_1), .COUTY1(na942_4), .IN1(~na1869_2), .IN2(na1063_2), .IN3(1'b1), .IN4(na1927_2), .IN5(1'b0), .IN6(1'b0),
                     .IN7(na1060_2), .IN8(na5_2), .CINX(1'b0), .CINY1(na941_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y75     80'h00_0018_00_0010_0666_80C4
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a943_1 ( .OUT(na943_1), .IN1(~na1869_2), .IN2(na1063_2), .IN3(1'b1), .IN4(na1929_2), .IN5(1'b0), .IN6(1'b0), .IN7(na2027_2),
                     .IN8(na5_2), .CINX(1'b0), .CINY1(na942_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y58     80'h00_0018_00_0010_0666_08A2
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a944_1 ( .OUT(na944_1), .COUTY1(na944_4), .IN1(na1225_1), .IN2(~na1054_1), .IN3(na1914_2), .IN4(1'b1), .IN5(na1061_2), .IN6(na1054_1),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na940_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y59     80'h00_0018_00_0010_0666_08C2
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a945_1 ( .OUT(na945_1), .COUTY1(na945_4), .IN1(na1226_2), .IN2(~na1054_1), .IN3(1'b1), .IN4(na250_1), .IN5(na1062_2), .IN6(na1054_1),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na944_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x93y60     80'h00_0078_00_0020_0C66_2C2C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a946_1 ( .OUT(na946_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na252_2), .IN7(na2040_2), .IN8(~na5_2),
                     .CINX(1'b0), .CINY1(na945_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a946_4 ( .OUT(na946_2), .COUTY1(na946_4), .IN1(1'b1), .IN2(na252_1), .IN3(na2039_2), .IN4(~na5_2), .IN5(1'b1), .IN6(na252_2),
                     .IN7(na2040_2), .IN8(~na5_2), .CINX(1'b0), .CINY1(na945_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x93y61     80'h00_0078_00_0020_0C66_2C2C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a948_1 ( .OUT(na948_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na254_2), .IN7(na2043_2), .IN8(~na5_2),
                     .CINX(1'b0), .CINY1(na946_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a948_4 ( .OUT(na948_2), .COUTY1(na948_4), .IN1(1'b1), .IN2(na254_1), .IN3(na2042_2), .IN4(~na5_2), .IN5(1'b1), .IN6(na254_2),
                     .IN7(na2043_2), .IN8(~na5_2), .CINX(1'b0), .CINY1(na946_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x93y62     80'h00_0078_00_0020_0C66_2C2C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a950_1 ( .OUT(na950_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na256_2), .IN7(na2045_2), .IN8(~na5_2),
                     .CINX(1'b0), .CINY1(na948_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a950_4 ( .OUT(na950_2), .COUTY1(na950_4), .IN1(1'b1), .IN2(na256_1), .IN3(na2044_2), .IN4(~na5_2), .IN5(1'b1), .IN6(na256_2),
                     .IN7(na2045_2), .IN8(~na5_2), .CINX(1'b0), .CINY1(na948_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y62     80'h00_0078_00_0020_0C66_A33A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a952_1 ( .OUT(na952_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na4_1), .IN7(na1496_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na1233_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a952_4 ( .OUT(na952_2), .COUTY1(na952_4), .IN1(na2103_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na7_1), .IN5(1'b1), .IN6(~na4_1),
                     .IN7(na1496_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na1233_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y67     80'h00_0078_00_0020_0C66_C3C3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a953_1 ( .OUT(na953_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na17_1), .IN7(1'b1), .IN8(na1463_1),
                     .CINX(1'b0), .CINY1(na982_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a953_4 ( .OUT(na953_2), .COUTY1(na953_4), .IN1(1'b1), .IN2(~na18_1), .IN3(1'b1), .IN4(na1459_2), .IN5(1'b1), .IN6(~na17_1),
                     .IN7(1'b1), .IN8(na1463_1), .CINX(1'b0), .CINY1(na982_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y68     80'h00_0078_00_0020_0C66_A5A3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a955_1 ( .OUT(na955_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na19_1), .IN6(1'b1), .IN7(na1455_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na953_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a955_4 ( .OUT(na955_2), .COUTY1(na955_4), .IN1(1'b1), .IN2(~na1886_2), .IN3(na1454_2), .IN4(1'b1), .IN5(~na19_1), .IN6(1'b1),
                     .IN7(na1455_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na953_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y69     80'h00_0078_00_0020_0C66_C5C5
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a957_1 ( .OUT(na957_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na21_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1452_1),
                     .CINX(1'b0), .CINY1(na955_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a957_4 ( .OUT(na957_2), .COUTY1(na957_4), .IN1(~na22_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1447_2), .IN5(~na21_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na1452_1), .CINX(1'b0), .CINY1(na955_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y70     80'h00_0078_00_0020_0C66_A5A3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a959_1 ( .OUT(na959_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na23_1), .IN6(1'b1), .IN7(na1442_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na957_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a959_4 ( .OUT(na959_2), .COUTY1(na959_4), .IN1(1'b1), .IN2(~na1888_2), .IN3(na1436_2), .IN4(1'b1), .IN5(~na23_1), .IN6(1'b1),
                     .IN7(na1442_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na957_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y71     80'h00_0078_00_0020_0C66_C3C3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a961_1 ( .OUT(na961_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na25_1), .IN7(1'b1), .IN8(na1433_1),
                     .CINX(1'b0), .CINY1(na959_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a961_4 ( .OUT(na961_2), .COUTY1(na961_4), .IN1(1'b1), .IN2(~na26_1), .IN3(1'b1), .IN4(na1430_2), .IN5(1'b1), .IN6(~na25_1),
                     .IN7(1'b1), .IN8(na1433_1), .CINX(1'b0), .CINY1(na959_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y72     80'h00_0078_00_0020_0C66_A5A3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a964_1 ( .OUT(na964_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na27_1), .IN6(1'b1), .IN7(na1525_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na961_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a964_4 ( .OUT(na964_2), .COUTY1(na964_4), .IN1(1'b1), .IN2(~na1891_2), .IN3(na1520_2), .IN4(1'b1), .IN5(~na27_1), .IN6(1'b1),
                     .IN7(na1525_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na961_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y73     80'h00_0078_00_0020_0C66_C5C3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a966_1 ( .OUT(na966_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na29_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1519_1),
                     .CINX(1'b0), .CINY1(na964_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a966_4 ( .OUT(na966_2), .COUTY1(na966_4), .IN1(1'b1), .IN2(~na30_1), .IN3(1'b1), .IN4(na1518_2), .IN5(~na29_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na1519_1), .CINX(1'b0), .CINY1(na964_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y74     80'h00_0078_00_0020_0C66_A3A5
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a968_1 ( .OUT(na968_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na1893_2), .IN7(na1517_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na966_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a968_4 ( .OUT(na968_2), .COUTY1(na968_4), .IN1(~na32_1), .IN2(1'b1), .IN3(na1516_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na1893_2),
                     .IN7(na1517_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na966_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y75     80'h00_0078_00_0020_0C66_C3C5
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a970_1 ( .OUT(na970_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na33_1), .IN7(1'b1), .IN8(na1514_1),
                     .CINX(1'b0), .CINY1(na968_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a970_4 ( .OUT(na970_2), .COUTY1(na970_4), .IN1(~na34_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1510_2), .IN5(1'b1), .IN6(~na33_1),
                     .IN7(1'b1), .IN8(na1514_1), .CINX(1'b0), .CINY1(na968_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y76     80'h00_0078_00_0020_0C66_A5A3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a972_1 ( .OUT(na972_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na35_1), .IN6(1'b1), .IN7(na1509_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na970_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a972_4 ( .OUT(na972_2), .COUTY1(na972_4), .IN1(1'b1), .IN2(~na1896_2), .IN3(na1504_2), .IN4(1'b1), .IN5(~na35_1), .IN6(1'b1),
                     .IN7(na1509_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na970_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y63     80'h00_0078_00_0020_0C66_C35C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a974_1 ( .OUT(na974_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na8_1), .IN7(1'b1), .IN8(na1492_1),
                     .CINX(1'b0), .CINY1(na952_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a974_4 ( .OUT(na974_2), .COUTY1(na974_4), .IN1(1'b1), .IN2(na2101_2), .IN3(~na10_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na8_1),
                     .IN7(1'b1), .IN8(na1492_1), .CINX(1'b0), .CINY1(na952_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y77     80'h00_0078_00_0020_0C66_C3C5
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a975_1 ( .OUT(na975_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na37_1), .IN7(1'b1), .IN8(na1503_1),
                     .CINX(1'b0), .CINY1(na972_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a975_4 ( .OUT(na975_2), .IN1(~na38_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1497_2), .IN5(1'b1), .IN6(~na37_1), .IN7(1'b1), .IN8(na1503_1),
                     .CINX(1'b0), .CINY1(na972_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y64     80'h00_0078_00_0020_0C66_3AA3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a978_1 ( .OUT(na978_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2100_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na11_1),
                     .CINX(1'b0), .CINY1(na974_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a978_4 ( .OUT(na978_2), .COUTY1(na978_4), .IN1(1'b1), .IN2(~na12_1), .IN3(na1480_2), .IN4(1'b1), .IN5(na2100_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(~na11_1), .CINX(1'b0), .CINY1(na974_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y65     80'h00_0078_00_0020_0C66_C3C5
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a980_1 ( .OUT(na980_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na13_1), .IN7(1'b1), .IN8(na1478_1),
                     .CINX(1'b0), .CINY1(na978_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a980_4 ( .OUT(na980_2), .COUTY1(na980_4), .IN1(~na14_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1475_2), .IN5(1'b1), .IN6(~na13_1),
                     .IN7(1'b1), .IN8(na1478_1), .CINX(1'b0), .CINY1(na978_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x75y66     80'h00_0078_00_0020_0C66_A5A3
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a982_1 ( .OUT(na982_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1881_2), .IN6(1'b1), .IN7(na1474_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na980_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a982_4 ( .OUT(na982_2), .COUTY1(na982_4), .IN1(1'b1), .IN2(~na16_1), .IN3(na1468_2), .IN4(1'b1), .IN5(~na1881_2), .IN6(1'b1),
                     .IN7(na1474_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na980_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y56     80'h00_0078_00_0020_0C66_ACCA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a984_1 ( .OUT(na984_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na4_1), .IN7(na1496_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na1239_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a984_4 ( .OUT(na984_2), .COUTY1(na984_4), .IN1(na2103_2), .IN2(1'b1), .IN3(1'b1), .IN4(na7_1), .IN5(1'b1), .IN6(na4_1), .IN7(na1496_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na1239_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y61     80'h00_0078_00_0020_0C66_CCCC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a985_1 ( .OUT(na985_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na17_1), .IN7(1'b1), .IN8(na1463_1),
                     .CINX(1'b0), .CINY1(na1015_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a985_4 ( .OUT(na985_2), .COUTY1(na985_4), .IN1(1'b1), .IN2(na18_1), .IN3(1'b1), .IN4(na1459_2), .IN5(1'b1), .IN6(na17_1),
                     .IN7(1'b1), .IN8(na1463_1), .CINX(1'b0), .CINY1(na1015_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y62     80'h00_0078_00_0020_0C66_AAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a987_1 ( .OUT(na987_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na19_1), .IN6(1'b1), .IN7(na1455_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na985_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a987_4 ( .OUT(na987_2), .COUTY1(na987_4), .IN1(1'b1), .IN2(na1886_2), .IN3(na1454_2), .IN4(1'b1), .IN5(na19_1), .IN6(1'b1),
                     .IN7(na1455_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na985_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y63     80'h00_0078_00_0020_0C66_CACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a989_1 ( .OUT(na989_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na21_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1452_1),
                     .CINX(1'b0), .CINY1(na987_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a989_4 ( .OUT(na989_2), .COUTY1(na989_4), .IN1(na22_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1447_2), .IN5(na21_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na1452_1), .CINX(1'b0), .CINY1(na987_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y64     80'h00_0078_00_0020_0C66_AAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a991_1 ( .OUT(na991_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na23_1), .IN6(1'b1), .IN7(na1442_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na989_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a991_4 ( .OUT(na991_2), .COUTY1(na991_4), .IN1(1'b1), .IN2(na1888_2), .IN3(na1436_2), .IN4(1'b1), .IN5(na23_1), .IN6(1'b1),
                     .IN7(na1442_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na989_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y65     80'h00_0078_00_0020_0C66_CCCC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a993_1 ( .OUT(na993_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na25_1), .IN7(1'b1), .IN8(na1433_1),
                     .CINX(1'b0), .CINY1(na991_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a993_4 ( .OUT(na993_2), .COUTY1(na993_4), .IN1(1'b1), .IN2(na26_1), .IN3(1'b1), .IN4(na1430_2), .IN5(1'b1), .IN6(na25_1),
                     .IN7(1'b1), .IN8(na1433_1), .CINX(1'b0), .CINY1(na991_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y66     80'h00_0078_00_0020_0C66_AAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a996_1 ( .OUT(na996_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na27_1), .IN6(1'b1), .IN7(na1525_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na993_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a996_4 ( .OUT(na996_2), .COUTY1(na996_4), .IN1(1'b1), .IN2(na1891_2), .IN3(na1520_2), .IN4(1'b1), .IN5(na27_1), .IN6(1'b1),
                     .IN7(na1525_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na993_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y67     80'h00_0078_00_0020_0C66_CACC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a998_1 ( .OUT(na998_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na29_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1519_1),
                     .CINX(1'b0), .CINY1(na996_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a998_4 ( .OUT(na998_2), .COUTY1(na998_4), .IN1(1'b1), .IN2(na30_1), .IN3(1'b1), .IN4(na1518_2), .IN5(na29_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na1519_1), .CINX(1'b0), .CINY1(na996_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y68     80'h00_0078_00_0020_0C66_ACAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1000_1 ( .OUT(na1000_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1893_2), .IN7(na1517_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na998_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1000_4 ( .OUT(na1000_2), .COUTY1(na1000_4), .IN1(na32_1), .IN2(1'b1), .IN3(na1516_2), .IN4(1'b1), .IN5(1'b1), .IN6(na1893_2),
                      .IN7(na1517_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na998_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y69     80'h00_0078_00_0020_0C66_CCCA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1002_1 ( .OUT(na1002_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na33_1), .IN7(1'b1), .IN8(na1514_1),
                      .CINX(1'b0), .CINY1(na1000_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1002_4 ( .OUT(na1002_2), .COUTY1(na1002_4), .IN1(na34_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1510_2), .IN5(1'b1), .IN6(na33_1),
                      .IN7(1'b1), .IN8(na1514_1), .CINX(1'b0), .CINY1(na1000_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y70     80'h00_0078_00_0020_0C66_AAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1004_1 ( .OUT(na1004_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na35_1), .IN6(1'b1), .IN7(na1509_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1002_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1004_4 ( .OUT(na1004_2), .COUTY1(na1004_4), .IN1(1'b1), .IN2(na1896_2), .IN3(na1504_2), .IN4(1'b1), .IN5(na35_1), .IN6(1'b1),
                      .IN7(na1509_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na1002_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y57     80'h00_0078_00_0020_0C66_CCAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1006_1 ( .OUT(na1006_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na8_1), .IN7(1'b1), .IN8(na1492_1),
                      .CINX(1'b0), .CINY1(na984_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1006_4 ( .OUT(na1006_2), .COUTY1(na1006_4), .IN1(1'b1), .IN2(na2101_2), .IN3(na10_1), .IN4(1'b1), .IN5(1'b1), .IN6(na8_1),
                      .IN7(1'b1), .IN8(na1492_1), .CINX(1'b0), .CINY1(na984_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y71     80'h00_0078_00_0020_0C66_CCCA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1007_1 ( .OUT(na1007_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na37_1), .IN7(1'b1), .IN8(na1503_1),
                      .CINX(1'b0), .CINY1(na1004_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1007_4 ( .OUT(na1007_2), .COUTY1(na1007_4), .IN1(na38_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1497_2), .IN5(1'b1), .IN6(na37_1),
                      .IN7(1'b1), .IN8(na1503_1), .CINX(1'b0), .CINY1(na1004_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x78y56     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1009_2 ( .OUT(na1009_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1009_6 ( .COUTY1(na1009_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1009_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x70y58     80'h00_0078_00_0020_0C66_CAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1011_1 ( .OUT(na1011_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2100_2), .IN6(1'b1), .IN7(1'b1), .IN8(na11_1),
                      .CINX(1'b0), .CINY1(na1006_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1011_4 ( .OUT(na1011_2), .COUTY1(na1011_4), .IN1(1'b1), .IN2(na12_1), .IN3(na1480_2), .IN4(1'b1), .IN5(na2100_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na11_1), .CINX(1'b0), .CINY1(na1006_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y59     80'h00_0078_00_0020_0C66_CCCA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1013_1 ( .OUT(na1013_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na13_1), .IN7(1'b1), .IN8(na1478_1),
                      .CINX(1'b0), .CINY1(na1011_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1013_4 ( .OUT(na1013_2), .COUTY1(na1013_4), .IN1(na14_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1475_2), .IN5(1'b1), .IN6(na13_1),
                      .IN7(1'b1), .IN8(na1478_1), .CINX(1'b0), .CINY1(na1011_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x70y60     80'h00_0078_00_0020_0C66_AAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1015_1 ( .OUT(na1015_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1881_2), .IN6(1'b1), .IN7(na1474_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1013_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1015_4 ( .OUT(na1015_2), .COUTY1(na1015_4), .IN1(1'b1), .IN2(na16_1), .IN3(na1468_2), .IN4(1'b1), .IN5(na1881_2), .IN6(1'b1),
                      .IN7(na1474_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na1013_4), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0000_0010)) 
           _a1018 ( .GLB0(na1018_1), .GLB1(_d3), .GLB2(_d4), .GLB3(_d5), .CLK_FB0(_d6), .CLK_FB1(_d7), .CLK_FB2(_d8), .CLK_FB3(_d9),
                    .CLK0_0(1'b0), .CLK0_90(1'b0), .CLK0_180(1'b0), .CLK0_270(1'b0), .CLK0_BYP(na40_1), .CLK1_0(1'b0), .CLK1_90(1'b0),
                    .CLK1_180(1'b0), .CLK1_270(1'b0), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0), .CLK2_270(1'b0),
                    .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0), .USR_GLB0(1'b0),
                    .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0), .USR_FB3(1'b0) );
// C_AND/D//AND/D      x87y56     80'h00_FE00_80_0000_0C88_AFF3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1023_1 ( .OUT(na1023_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na862_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1023_2 ( .OUT(na1023_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1023_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1023_4 ( .OUT(na1023_2_i), .IN1(1'b1), .IN2(~na1023_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1023_5 ( .OUT(na1023_2), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1023_2_i) );
// C_AND/D///      x93y54     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1025_1 ( .OUT(na1025_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na876_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1025_2 ( .OUT(na1025_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1025_1_i) );
// C_///AND/D      x92y56     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1027_4 ( .OUT(na1027_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na878_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1027_5 ( .OUT(na1027_2), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1027_2_i) );
// C_AND/D///      x91y55     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1029_1 ( .OUT(na1029_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na880_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1029_2 ( .OUT(na1029_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1029_1_i) );
// C_///AND/D      x91y57     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1031_4 ( .OUT(na1031_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na882_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1031_5 ( .OUT(na1031_2), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1031_2_i) );
// C_///AND/D      x89y59     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1033_4 ( .OUT(na1033_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na853_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1033_5 ( .OUT(na1033_2), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1033_2_i) );
// C_AND/D///      x91y58     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1035_1 ( .OUT(na1035_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na855_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1035_2 ( .OUT(na1035_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1035_1_i) );
// C_AND/D///      x91y59     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1037_1 ( .OUT(na1037_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na857_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1037_2 ( .OUT(na1037_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1037_1_i) );
// C_AND/D///      x94y61     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1039_1 ( .OUT(na1039_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na859_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1039_2 ( .OUT(na1039_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1039_1_i) );
// C_///AND/D      x91y59     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1041_4 ( .OUT(na1041_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na861_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1041_5 ( .OUT(na1041_2), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1041_2_i) );
// C_AND/D///      x94y60     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1043_1 ( .OUT(na1043_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na864_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1043_2 ( .OUT(na1043_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1043_1_i) );
// C_///AND/D      x88y61     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1045_4 ( .OUT(na1045_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na866_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1045_5 ( .OUT(na1045_2), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1045_2_i) );
// C_///AND/D      x88y63     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1047_4 ( .OUT(na1047_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na868_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1047_5 ( .OUT(na1047_2), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1047_2_i) );
// C_///AND/D      x94y65     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1049_4 ( .OUT(na1049_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na870_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1049_5 ( .OUT(na1049_2), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1049_2_i) );
// C_AND/D///      x88y61     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1051_1 ( .OUT(na1051_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na872_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1051_2 ( .OUT(na1051_1), .CLK(na1018_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1051_1_i) );
// C_///AND/D      x85y63     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1053_4 ( .OUT(na1053_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1154_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1053_5 ( .OUT(na1053_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1053_2_i) );
// C_AND/D///      x89y58     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1054_1 ( .OUT(na1054_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1165_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1054_2 ( .OUT(na1054_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1054_1_i) );
// C_AND/D//AND/D      x86y61     80'h00_FA00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1055_1 ( .OUT(na1055_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1168_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1055_2 ( .OUT(na1055_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1055_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1055_4 ( .OUT(na1055_2_i), .IN1(na1170_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1055_5 ( .OUT(na1055_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1055_2_i) );
// C_AND/D///      x82y58     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1056_1 ( .OUT(na1056_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1169_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1056_2 ( .OUT(na1056_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1056_1_i) );
// C_AND/D//AND/D      x81y53     80'h00_FA00_80_0000_0C88_FCCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1058_1 ( .OUT(na1058_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1171_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1058_2 ( .OUT(na1058_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1058_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1058_4 ( .OUT(na1058_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1155_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1058_5 ( .OUT(na1058_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1058_2_i) );
// C_AND/D//AND/D      x77y53     80'h00_FA00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1059_1 ( .OUT(na1059_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1172_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1059_2 ( .OUT(na1059_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1059_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1059_4 ( .OUT(na1059_2_i), .IN1(na1156_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1059_5 ( .OUT(na1059_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1059_2_i) );
// C_AND/D//AND/D      x80y57     80'h00_FA00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1060_1 ( .OUT(na1060_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1173_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1060_2 ( .OUT(na1060_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1060_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1060_4 ( .OUT(na1060_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1157_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1060_5 ( .OUT(na1060_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1060_2_i) );
// C_AND/D//AND/D      x81y59     80'h00_FA00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1061_1 ( .OUT(na1061_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1144_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1061_2 ( .OUT(na1061_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1061_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1061_4 ( .OUT(na1061_2_i), .IN1(na1158_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1061_5 ( .OUT(na1061_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1061_2_i) );
// C_AND/D//AND/D      x79y55     80'h00_FA00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1062_1 ( .OUT(na1062_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1062_2 ( .OUT(na1062_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1062_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1062_4 ( .OUT(na1062_2_i), .IN1(na1159_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1062_5 ( .OUT(na1062_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1062_2_i) );
// C_AND/D//AND/D      x77y58     80'h00_FA00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1063_1 ( .OUT(na1063_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1063_2 ( .OUT(na1063_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1063_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1063_4 ( .OUT(na1063_2_i), .IN1(na1167_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1063_5 ( .OUT(na1063_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1063_2_i) );
// C_AND/D///      x81y57     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1064_1 ( .OUT(na1064_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1064_2 ( .OUT(na1064_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1064_1_i) );
// C_///AND/D      x82y60     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1065_4 ( .OUT(na1065_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1148_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1065_5 ( .OUT(na1065_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1065_2_i) );
// C_AND/D///      x90y66     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1066_1 ( .OUT(na1066_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1149_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1066_2 ( .OUT(na1066_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1066_1_i) );
// C_///AND/D      x90y66     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1067_4 ( .OUT(na1067_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1150_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1067_5 ( .OUT(na1067_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1067_2_i) );
// C_///AND/D      x92y66     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1068_4 ( .OUT(na1068_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1151_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1068_5 ( .OUT(na1068_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1068_2_i) );
// C_///AND/D      x90y68     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1069_4 ( .OUT(na1069_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1152_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1069_5 ( .OUT(na1069_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1069_2_i) );
// C_AND/D///      x92y68     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1070_1 ( .OUT(na1070_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1153_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1070_2 ( .OUT(na1070_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1070_1_i) );
// C_AND/D//AND/D      x81y55     80'h00_FA00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1077_1 ( .OUT(na1077_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1161_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1077_2 ( .OUT(na1077_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1077_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1077_4 ( .OUT(na1077_2_i), .IN1(na1160_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1077_5 ( .OUT(na1077_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1077_2_i) );
// C_AND/D//AND/D      x83y59     80'h00_FA00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1079_1 ( .OUT(na1079_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1163_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1079_2 ( .OUT(na1079_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1079_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1079_4 ( .OUT(na1079_2_i), .IN1(na1162_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1079_5 ( .OUT(na1079_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1079_2_i) );
// C_AND/D//AND/D      x83y53     80'h00_FA00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1081_1 ( .OUT(na1081_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1166_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1081_2 ( .OUT(na1081_1), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1081_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1081_4 ( .OUT(na1081_2_i), .IN1(na1164_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1081_5 ( .OUT(na1081_2), .CLK(na1018_1), .EN(na240_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1081_2_i) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a1108 ( .Y(na1108_1), .I(clk) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1109 ( .O(mem_addr[0]), .A(na1797_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1110 ( .O(mem_addr[1]), .A(na1798_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1111 ( .O(mem_addr[10]), .A(na1799_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1112 ( .O(mem_addr[11]), .A(na1800_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1113 ( .O(mem_addr[12]), .A(na1801_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1114 ( .O(mem_addr[13]), .A(na1802_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1115 ( .O(mem_addr[14]), .A(na1803_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1116 ( .O(mem_addr[15]), .A(na1804_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1117 ( .O(mem_addr[16]), .A(na1805_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1118 ( .O(mem_addr[17]), .A(na1806_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1119 ( .O(mem_addr[18]), .A(na1807_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1120 ( .O(mem_addr[19]), .A(na1808_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1121 ( .O(mem_addr[2]), .A(na1809_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1122 ( .O(mem_addr[20]), .A(na1810_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1123 ( .O(mem_addr[21]), .A(na1811_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1124 ( .O(mem_addr[22]), .A(na1812_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1125 ( .O(mem_addr[23]), .A(na1813_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1126 ( .O(mem_addr[24]), .A(na1814_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1127 ( .O(mem_addr[25]), .A(na1815_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1128 ( .O(mem_addr[26]), .A(na1816_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1129 ( .O(mem_addr[27]), .A(na1817_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1130 ( .O(mem_addr[28]), .A(na1818_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1131 ( .O(mem_addr[29]), .A(na1819_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1132 ( .O(mem_addr[3]), .A(na1820_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1133 ( .O(mem_addr[30]), .A(na1821_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1134 ( .O(mem_addr[31]), .A(na1822_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1135 ( .O(mem_addr[4]), .A(na1823_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1136 ( .O(mem_addr[5]), .A(na1824_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1137 ( .O(mem_addr[6]), .A(na1825_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1138 ( .O(mem_addr[7]), .A(na1826_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1139 ( .O(mem_addr[8]), .A(na1827_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1140 ( .O(mem_addr[9]), .A(na1828_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1141 ( .Y(na1141_1), .I(mem_rbusy) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1142 ( .Y(na1142_1), .I(mem_rdata[0]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1143 ( .Y(na1143_1), .I(mem_rdata[1]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1144 ( .Y(na1144_1), .I(mem_rdata[10]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1145 ( .Y(na1145_1), .I(mem_rdata[11]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1146 ( .Y(na1146_1), .I(mem_rdata[12]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1147 ( .Y(na1147_1), .I(mem_rdata[13]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1148 ( .Y(na1148_1), .I(mem_rdata[14]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1149 ( .Y(na1149_1), .I(mem_rdata[15]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1150 ( .Y(na1150_1), .I(mem_rdata[16]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1151 ( .Y(na1151_1), .I(mem_rdata[17]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1152 ( .Y(na1152_1), .I(mem_rdata[18]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1153 ( .Y(na1153_1), .I(mem_rdata[19]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1154 ( .Y(na1154_1), .I(mem_rdata[2]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1155 ( .Y(na1155_1), .I(mem_rdata[20]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1156 ( .Y(na1156_1), .I(mem_rdata[21]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1157 ( .Y(na1157_1), .I(mem_rdata[22]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1158 ( .Y(na1158_1), .I(mem_rdata[23]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1159 ( .Y(na1159_1), .I(mem_rdata[24]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1160 ( .Y(na1160_1), .I(mem_rdata[25]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1161 ( .Y(na1161_1), .I(mem_rdata[26]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1162 ( .Y(na1162_1), .I(mem_rdata[27]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1163 ( .Y(na1163_1), .I(mem_rdata[28]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1164 ( .Y(na1164_1), .I(mem_rdata[29]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1165 ( .Y(na1165_1), .I(mem_rdata[3]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1166 ( .Y(na1166_1), .I(mem_rdata[30]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1167 ( .Y(na1167_1), .I(mem_rdata[31]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1168 ( .Y(na1168_1), .I(mem_rdata[4]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1169 ( .Y(na1169_1), .I(mem_rdata[5]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1170 ( .Y(na1170_1), .I(mem_rdata[6]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1171 ( .Y(na1171_1), .I(mem_rdata[7]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1172 ( .Y(na1172_1), .I(mem_rdata[8]) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1173 ( .Y(na1173_1), .I(mem_rdata[9]) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1174 ( .O(mem_rstrb), .A(na1829_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1175 ( .Y(na1175_1), .I(mem_wbusy) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1176 ( .O(mem_wdata[0]), .A(na1830_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1177 ( .O(mem_wdata[1]), .A(na1831_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1178 ( .O(mem_wdata[10]), .A(na1832_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1179 ( .O(mem_wdata[11]), .A(na1833_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1180 ( .O(mem_wdata[12]), .A(na1834_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1181 ( .O(mem_wdata[13]), .A(na1835_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1182 ( .O(mem_wdata[14]), .A(na1836_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1183 ( .O(mem_wdata[15]), .A(na1837_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1184 ( .O(mem_wdata[16]), .A(na1838_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1185 ( .O(mem_wdata[17]), .A(na1839_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1186 ( .O(mem_wdata[18]), .A(na1840_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1187 ( .O(mem_wdata[19]), .A(na1841_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1188 ( .O(mem_wdata[2]), .A(na1842_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1189 ( .O(mem_wdata[20]), .A(na1843_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1190 ( .O(mem_wdata[21]), .A(na1844_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1191 ( .O(mem_wdata[22]), .A(na1845_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1192 ( .O(mem_wdata[23]), .A(na1846_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1193 ( .O(mem_wdata[24]), .A(na1847_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1194 ( .O(mem_wdata[25]), .A(na1848_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1195 ( .O(mem_wdata[26]), .A(na1849_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1196 ( .O(mem_wdata[27]), .A(na1850_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1197 ( .O(mem_wdata[28]), .A(na1851_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1198 ( .O(mem_wdata[29]), .A(na1852_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1199 ( .O(mem_wdata[3]), .A(na1853_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1200 ( .O(mem_wdata[30]), .A(na1854_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1201 ( .O(mem_wdata[31]), .A(na1855_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1202 ( .O(mem_wdata[4]), .A(na1856_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1203 ( .O(mem_wdata[5]), .A(na1857_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1204 ( .O(mem_wdata[6]), .A(na1858_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1205 ( .O(mem_wdata[7]), .A(na1859_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1206 ( .O(mem_wdata[8]), .A(na1860_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1207 ( .O(mem_wdata[9]), .A(na1861_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1208 ( .O(mem_wmask[0]), .A(na1862_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1209 ( .O(mem_wmask[1]), .A(na1863_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1210 ( .O(mem_wmask[2]), .A(na1864_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1211 ( .O(mem_wmask[3]), .A(na1865_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000050)) 
           _a1212 ( .Y(na1212_1), .I(reset) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_00_06_00_00_C3_03_00_23_00_00_23_00_13_23_00_00_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a1213 ( .DOA({na1213_1, na1213_2, na1213_3, na1213_4, na1213_5, na1213_6, na1213_7, na1213_8, na1213_9, na1213_10, na1213_11,
                   na1213_12, na1213_13, na1213_14, na1213_15, na1213_16, na1213_17, na1213_18, na1213_19, na1213_20, _d10, _d11, _d12,
                   _d13, _d14, _d15, _d16, _d17, _d18, _d19, _d20, _d21, _d22, _d23, _d24, _d25, _d26, _d27, _d28, _d29}),
                    .DOAX({_d30, _d31, _d32, _d33, _d34, _d35, _d36, _d37, _d38, _d39, _d40, _d41, _d42, _d43, _d44, _d45, _d46, _d47,
                   _d48, _d49, _d50, _d51, _d52, _d53, _d54, _d55, _d56, _d57, _d58, _d59, _d60, _d61, _d62, _d63, _d64, _d65, _d66,
                   _d67, _d68, _d69}),
                    .DOB({_d70, _d71, _d72, _d73, _d74, _d75, _d76, _d77, na1213_89, na1213_90, na1213_91, na1213_92, na1213_93, na1213_94,
                   na1213_95, na1213_96, na1213_97, na1213_98, na1213_99, na1213_100, _d78, _d79, _d80, _d81, _d82, _d83, _d84, _d85,
                   _d86, _d87, _d88, _d89, _d90, _d91, _d92, _d93, _d94, _d95, _d96, _d97}),
                    .DOBX({_d98, _d99, _d100, _d101, _d102, _d103, _d104, _d105, _d106, _d107, _d108, _d109, _d110, _d111, _d112, _d113,
                   _d114, _d115, _d116, _d117, _d118, _d119, _d120, _d121, _d122, _d123, _d124, _d125, _d126, _d127, _d128, _d129, _d130,
                   _d131, _d132, _d133, _d134, _d135, _d136, _d137}),
                    .ECC1B_ERRA({_d138, _d139, _d140, _d141}),
                    .ECC1B_ERRB({_d142, _d143, _d144, _d145}),
                    .ECC2B_ERRA({_d146, _d147, _d148, _d149}),
                    .ECC2B_ERRB({_d150, _d151, _d152, _d153}),
                    .FORW_CAS_WRAO(_d154), .FORW_CAS_WRBO(_d155), .FORW_CAS_BMAO(_d156), .FORW_CAS_BMBO(_d157), .FORW_CAS_RDAO(_d158),
                    .FORW_CAS_RDBO(_d159), .FORW_UADDRAO({_d160, _d161, _d162, _d163, _d164, _d165, _d166, _d167, _d168, _d169, _d170,
                   _d171, _d172, _d173, _d174, _d175}),
                    .FORW_LADDRAO({_d176, _d177, _d178, _d179, _d180, _d181, _d182, _d183, _d184, _d185, _d186, _d187, _d188, _d189,
                   _d190, _d191}),
                    .FORW_UADDRBO({_d192, _d193, _d194, _d195, _d196, _d197, _d198, _d199, _d200, _d201, _d202, _d203, _d204, _d205,
                   _d206, _d207}),
                    .FORW_LADDRBO({_d208, _d209, _d210, _d211, _d212, _d213, _d214, _d215, _d216, _d217, _d218, _d219, _d220, _d221,
                   _d222, _d223}),
                    .FORW_UA0CLKO(_d224), .FORW_UA0ENO(_d225), .FORW_UA0WEO(_d226), .FORW_LA0CLKO(_d227), .FORW_LA0ENO(_d228), .FORW_LA0WEO(_d229),
                    .FORW_UA1CLKO(_d230), .FORW_UA1ENO(_d231), .FORW_UA1WEO(_d232), .FORW_LA1CLKO(_d233), .FORW_LA1ENO(_d234), .FORW_LA1WEO(_d235),
                    .FORW_UB0CLKO(_d236), .FORW_UB0ENO(_d237), .FORW_UB0WEO(_d238), .FORW_LB0CLKO(_d239), .FORW_LB0ENO(_d240), .FORW_LB0WEO(_d241),
                    .FORW_UB1CLKO(_d242), .FORW_UB1ENO(_d243), .FORW_UB1WEO(_d244), .FORW_LB1CLKO(_d245), .FORW_LB1ENO(_d246), .FORW_LB1WEO(_d247),
                    .CLOCKA({_d248, _d249, _d250, _d251}),
                    .CLOCKB({_d252, _d253, _d254, _d255}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, na1215_9, 1'b1, 1'b1}),
                    .GLWEA({1'b1, na1217_10, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1({na1219_10, na1221_9, na1230_10, na1234_9, na1237_10, na1238_9, na1241_10, na1242_9, na1245_10, na1246_9,
                   na1247_10, na1249_9, na1250_10, na1251_9, na1253_10, na1254_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({na1255_10, na1257_9, na1258_10, na1259_9, na1261_10, na1262_9, na1263_10, na1265_9, na1266_10, na1267_9,
                   na1269_10, na1270_9, na1271_10, na1273_9, na1274_10, na1275_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na1277_10, na1278_9, na1279_10, na1281_9, na1282_10, na1283_9, na1285_10, na1286_9, na1287_10, na1289_9, na1290_10,
                   na1291_9, na1293_10, na1294_9, na1295_10, na1297_9, na1298_10, na1299_9, na1301_10, na1302_9, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na1303_10, na1305_9, na1306_10, na1307_9, na1309_10, na1310_9,
                   na1311_10, na1313_9, na1314_10, na1315_9, na1317_10, na1318_9, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({na1319_10, na1321_9, na1322_10, na1323_9, na1324_10, na1325_9, na1328_10, na1330_9, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na1018_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_00_00_C0_00_1B_00_00_23_03_00_23_00_00_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a1214 ( .DOA({_d256, _d257, _d258, _d259, _d260, _d261, _d262, _d263, _d264, _d265, _d266, _d267, _d268, _d269, _d270, _d271,
                   _d272, _d273, _d274, _d275, na1214_21, na1214_22, na1214_23, na1214_24, na1214_25, na1214_26, na1214_27, na1214_28,
                   na1214_29, na1214_30, na1214_31, na1214_32, na1214_33, na1214_34, na1214_35, na1214_36, na1214_37, na1214_38, na1214_39,
                   na1214_40}),
                    .DOAX({_d276, _d277, _d278, _d279, _d280, _d281, _d282, _d283, _d284, _d285, _d286, _d287, _d288, _d289, _d290,
                   _d291, _d292, _d293, _d294, _d295, _d296, _d297, _d298, _d299, _d300, _d301, _d302, _d303, _d304, _d305, _d306, _d307,
                   _d308, _d309, _d310, _d311, _d312, _d313, _d314, _d315}),
                    .DOB({_d316, _d317, _d318, _d319, _d320, _d321, _d322, _d323, _d324, _d325, _d326, _d327, _d328, _d329, _d330, _d331,
                   _d332, _d333, _d334, _d335, _d336, _d337, _d338, _d339, _d340, _d341, _d342, _d343, na1214_109, na1214_110, na1214_111,
                   na1214_112, na1214_113, na1214_114, na1214_115, na1214_116, na1214_117, na1214_118, na1214_119, na1214_120}),
                    .DOBX({_d344, _d345, _d346, _d347, _d348, _d349, _d350, _d351, _d352, _d353, _d354, _d355, _d356, _d357, _d358,
                   _d359, _d360, _d361, _d362, _d363, _d364, _d365, _d366, _d367, _d368, _d369, _d370, _d371, _d372, _d373, _d374, _d375,
                   _d376, _d377, _d378, _d379, _d380, _d381, _d382, _d383}),
                    .ECC1B_ERRA({_d384, _d385, _d386, _d387}),
                    .ECC1B_ERRB({_d388, _d389, _d390, _d391}),
                    .ECC2B_ERRA({_d392, _d393, _d394, _d395}),
                    .ECC2B_ERRB({_d396, _d397, _d398, _d399}),
                    .FORW_CAS_WRAO(_d400), .FORW_CAS_WRBO(_d401), .FORW_CAS_BMAO(_d402), .FORW_CAS_BMBO(_d403), .FORW_CAS_RDAO(_d404),
                    .FORW_CAS_RDBO(_d405), .FORW_UADDRAO({_d406, _d407, _d408, _d409, _d410, _d411, _d412, _d413, _d414, _d415, _d416,
                   _d417, _d418, _d419, _d420, _d421}),
                    .FORW_LADDRAO({_d422, _d423, _d424, _d425, _d426, _d427, _d428, _d429, _d430, _d431, _d432, _d433, _d434, _d435,
                   _d436, _d437}),
                    .FORW_UADDRBO({_d438, _d439, _d440, _d441, _d442, _d443, _d444, _d445, _d446, _d447, _d448, _d449, _d450, _d451,
                   _d452, _d453}),
                    .FORW_LADDRBO({_d454, _d455, _d456, _d457, _d458, _d459, _d460, _d461, _d462, _d463, _d464, _d465, _d466, _d467,
                   _d468, _d469}),
                    .FORW_UA0CLKO(_d470), .FORW_UA0ENO(_d471), .FORW_UA0WEO(_d472), .FORW_LA0CLKO(_d473), .FORW_LA0ENO(_d474), .FORW_LA0WEO(_d475),
                    .FORW_UA1CLKO(_d476), .FORW_UA1ENO(_d477), .FORW_UA1WEO(_d478), .FORW_LA1CLKO(_d479), .FORW_LA1ENO(_d480), .FORW_LA1WEO(_d481),
                    .FORW_UB0CLKO(_d482), .FORW_UB0ENO(_d483), .FORW_UB0WEO(_d484), .FORW_LB0CLKO(_d485), .FORW_LB0ENO(_d486), .FORW_LB0WEO(_d487),
                    .FORW_UB1CLKO(_d488), .FORW_UB1ENO(_d489), .FORW_UB1WEO(_d490), .FORW_LB1CLKO(_d491), .FORW_LB1ENO(_d492), .FORW_LB1WEO(_d493),
                    .CLOCKA({_d494, _d495, _d496, _d497}),
                    .CLOCKB({_d498, _d499, _d500, _d501}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, na1334_9}),
                    .GLWEA({1'b1, 1'b1, 1'b1, na1335_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na1338_10, na1339_9, na1340_10, na1343_9, na1344_10, na1345_9, na1354_10, na1358_9, na1360_10, na1363_9,
                   na1367_10, na1368_9, na1369_10, na1371_9, na1373_10, na1378_9}),
                    .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({na1380_10, na1381_9, na1385_10, na1387_9, na1388_10, na1392_9, na1398_10, na1403_9, na1404_10, na1405_9,
                   na1406_10, na1409_9, na1416_10, na1419_9, na1423_10, na1425_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, na1430_10, na1433_9, na1436_10, na1442_9, na1447_10, na1452_9, na1454_10, na1455_9, na1459_10, na1463_9,
                   na1468_10, na1474_9, na1475_10, na1478_9, na1480_10, na1484_9, na1491_10, na1492_9, na1493_10, na1496_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na1497_10, na1503_9, na1504_10, na1509_9, na1510_10,
                   na1514_9, na1516_10, na1517_9, na1518_10, na1519_9, na1520_10, na1525_9}),
                    .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, na1526_10, na1530_9, na1533_10, na1534_9, na1535_10, na1539_9, na1540_10, na1546_9, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na1018_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
// C_AND////      x67y58     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1215_1 ( .OUT(na1215_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na240_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1215_6 ( .RAM_O1(na1215_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1215_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x88y72     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1216_4 ( .OUT(na1216_2), .IN1(na1141_1), .IN2(1'b1), .IN3(na42_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x59y57     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1217_4 ( .OUT(na1217_2), .IN1(1'b1), .IN2(na39_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1217_6 ( .RAM_O2(na1217_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1217_2), .COMP_OUT(1'b0) );
// C_///AND/      x86y71     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1218_4 ( .OUT(na1218_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na240_2), .IN4(~na241_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1219_4 ( .OUT(na1219_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1219_6 ( .RAM_O2(na1219_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1219_2), .COMP_OUT(1'b0) );
// C_AND////      x79y51     80'h00_0018_00_0000_0888_F151
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1220_1 ( .OUT(na1220_1), .IN1(~na1059_1), .IN2(~na2022_2), .IN3(~na1060_1), .IN4(1'b1), .IN5(~na1062_1), .IN6(~na2026_2),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1221_1 ( .OUT(na1221_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1221_6 ( .RAM_O1(na1221_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1221_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x95y61     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1222_2 ( .OUT(na1222_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1222_6 ( .COUTY1(na1222_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1222_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x83y61     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1223_4 ( .OUT(na1223_2), .IN1(na1059_1), .IN2(1'b1), .IN3(~na1055_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x83y57     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1224_1 ( .OUT(na1224_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2019_2), .IN6(1'b1), .IN7(na1060_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y53     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1225_1 ( .OUT(na1225_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1061_1), .IN6(1'b1), .IN7(~na1055_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y61     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1226_4 ( .OUT(na1226_2), .IN1(na1062_1), .IN2(1'b1), .IN3(~na1055_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y63     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1227_4 ( .OUT(na1227_2), .IN1(na1058_1), .IN2(1'b1), .IN3(~na1055_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x87y76     80'h00_0078_00_0000_0C88_3A2F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1228_1 ( .OUT(na1228_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na47_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na44_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1228_4 ( .OUT(na1228_2), .IN1(1'b1), .IN2(1'b1), .IN3(na240_2), .IN4(~na44_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x80y75     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1229_1 ( .OUT(na1229_1), .IN1(~na78_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1981_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1230_4 ( .OUT(na1230_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1230_6 ( .RAM_O2(na1230_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1230_2), .COMP_OUT(1'b0) );
// C_AND////      x89y68     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1231_1 ( .OUT(na1231_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na86_1), .IN7(1'b1), .IN8(na81_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x93y55     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1232_2 ( .OUT(na1232_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1232_6 ( .COUTY1(na1232_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1232_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x75y61     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1233_2 ( .OUT(na1233_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1233_6 ( .COUTY1(na1233_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1233_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x60y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1234_1 ( .OUT(na1234_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1234_6 ( .RAM_O1(na1234_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1234_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x93y81     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1235_4 ( .OUT(na1235_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na42_1), .IN4(~na50_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x82y78     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1236_1 ( .OUT(na1236_1), .IN1(~na107_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1986_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y62     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1237_4 ( .OUT(na1237_2), .IN1(na1062_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1237_6 ( .RAM_O2(na1237_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1237_2), .COMP_OUT(1'b0) );
// C_AND////      x60y62     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1238_1 ( .OUT(na1238_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1061_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1238_6 ( .RAM_O1(na1238_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1238_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x70y55     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1239_2 ( .OUT(na1239_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1239_6 ( .COUTY1(na1239_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1239_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x94y74     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1240_1 ( .OUT(na1240_1), .IN1(~na112_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1987_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y61     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1241_4 ( .OUT(na1241_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1060_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1241_6 ( .RAM_O2(na1241_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1241_2), .COMP_OUT(1'b0) );
// C_AND////      x60y61     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1242_1 ( .OUT(na1242_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1059_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1242_6 ( .RAM_O1(na1242_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1242_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x70y72     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a1243_1 ( .OUT(na1243_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1007_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x96y72     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1244_1 ( .OUT(na1244_1), .IN1(~na117_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1988_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y60     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1245_4 ( .OUT(na1245_2), .IN1(na1058_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1245_6 ( .RAM_O2(na1245_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1245_2), .COMP_OUT(1'b0) );
// C_AND////      x60y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1246_1 ( .OUT(na1246_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1246_6 ( .RAM_O1(na1246_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1246_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y59     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1247_4 ( .OUT(na1247_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1247_6 ( .RAM_O2(na1247_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1247_2), .COMP_OUT(1'b0) );
// C_ORAND////      x98y75     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1248_1 ( .OUT(na1248_1), .IN1(~na122_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1989_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y59     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1249_1 ( .OUT(na1249_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1249_6 ( .RAM_O1(na1249_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1249_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y58     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1250_4 ( .OUT(na1250_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1250_6 ( .RAM_O2(na1250_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1250_2), .COMP_OUT(1'b0) );
// C_AND////      x60y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1251_1 ( .OUT(na1251_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1251_6 ( .RAM_O1(na1251_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1251_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x100y71     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1252_1 ( .OUT(na1252_1), .IN1(~na127_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1990_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1253_4 ( .OUT(na1253_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1253_6 ( .RAM_O2(na1253_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1253_2), .COMP_OUT(1'b0) );
// C_AND////      x60y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1254_1 ( .OUT(na1254_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1254_6 ( .RAM_O1(na1254_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1254_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1255_4 ( .OUT(na1255_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1255_6 ( .RAM_O2(na1255_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1255_2), .COMP_OUT(1'b0) );
// C_ORAND////      x100y73     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1256_1 ( .OUT(na1256_1), .IN1(~na132_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1991_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1257_1 ( .OUT(na1257_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1257_6 ( .RAM_O1(na1257_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1257_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1258_4 ( .OUT(na1258_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1258_6 ( .RAM_O2(na1258_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1258_2), .COMP_OUT(1'b0) );
// C_AND////      x69y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1259_1 ( .OUT(na1259_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1259_6 ( .RAM_O1(na1259_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1259_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x100y74     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1260_1 ( .OUT(na1260_1), .IN1(~na137_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1992_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y62     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1261_4 ( .OUT(na1261_2), .IN1(na1159_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1261_6 ( .RAM_O2(na1261_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1261_2), .COMP_OUT(1'b0) );
// C_AND////      x69y62     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1262_1 ( .OUT(na1262_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1158_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1262_6 ( .RAM_O1(na1262_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1262_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y61     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1263_4 ( .OUT(na1263_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1157_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1263_6 ( .RAM_O2(na1263_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1263_2), .COMP_OUT(1'b0) );
// C_ORAND////      x96y74     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1264_1 ( .OUT(na1264_1), .IN1(~na142_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1993_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y61     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1265_1 ( .OUT(na1265_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1156_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1265_6 ( .RAM_O1(na1265_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1265_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y60     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1266_4 ( .OUT(na1266_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1155_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1266_6 ( .RAM_O2(na1266_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1266_2), .COMP_OUT(1'b0) );
// C_AND////      x69y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1267_1 ( .OUT(na1267_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1267_6 ( .RAM_O1(na1267_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1267_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x92y76     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1268_1 ( .OUT(na1268_1), .IN1(~na147_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1994_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y59     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1269_4 ( .OUT(na1269_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1269_6 ( .RAM_O2(na1269_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1269_2), .COMP_OUT(1'b0) );
// C_AND////      x69y59     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1270_1 ( .OUT(na1270_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1270_6 ( .RAM_O1(na1270_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1270_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y58     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1271_4 ( .OUT(na1271_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1271_6 ( .RAM_O2(na1271_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1271_2), .COMP_OUT(1'b0) );
// C_ORAND////      x80y79     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1272_1 ( .OUT(na1272_1), .IN1(~na152_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1971_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1273_1 ( .OUT(na1273_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1273_6 ( .RAM_O1(na1273_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1273_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1274_4 ( .OUT(na1274_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1274_6 ( .RAM_O2(na1274_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1274_2), .COMP_OUT(1'b0) );
// C_AND////      x69y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1275_1 ( .OUT(na1275_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1275_6 ( .RAM_O1(na1275_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1275_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x84y79     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1276_1 ( .OUT(na1276_1), .IN1(~na157_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1972_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x62y64     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1277_4 ( .OUT(na1277_2_i), .IN1(na827_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1277_5 ( .OUT(na1277_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_1), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1277_6 ( .RAM_O2(na1277_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1277_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x62y64     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1278_1 ( .OUT(na1278_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na824_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1278_2 ( .OUT(na1278_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_2), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1278_6 ( .RAM_O1(na1278_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1278_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x62y63     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1279_4 ( .OUT(na1279_2_i), .IN1(1'b1), .IN2(na616_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1279_5 ( .OUT(na1279_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_3), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1279_6 ( .RAM_O2(na1279_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1279_2_i), .COMP_OUT(1'b0) );
// C_ORAND////      x86y77     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1280_1 ( .OUT(na1280_1), .IN1(~na162_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1973_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x62y63     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1281_1 ( .OUT(na1281_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na821_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1281_2 ( .OUT(na1281_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_4), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1281_6 ( .RAM_O1(na1281_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1281_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y64     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1282_4 ( .OUT(na1282_2_i), .IN1(1'b1), .IN2(na594_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1282_5 ( .OUT(na1282_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_5), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1282_6 ( .RAM_O2(na1282_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1282_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y64     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1283_1 ( .OUT(na1283_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na581_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1283_2 ( .OUT(na1283_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_6), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1283_6 ( .RAM_O1(na1283_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1283_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x90y77     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1284_1 ( .OUT(na1284_1), .IN1(~na167_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1974_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y63     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1285_4 ( .OUT(na1285_2_i), .IN1(na568_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1285_5 ( .OUT(na1285_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_7), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1285_6 ( .RAM_O2(na1285_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1285_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y63     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1286_1 ( .OUT(na1286_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na812_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1286_2 ( .OUT(na1286_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_8), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1286_6 ( .RAM_O1(na1286_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1286_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y62     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1287_4 ( .OUT(na1287_2_i), .IN1(na809_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1287_5 ( .OUT(na1287_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_9), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1287_6 ( .RAM_O2(na1287_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1287_2_i), .COMP_OUT(1'b0) );
// C_ORAND////      x90y83     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1288_1 ( .OUT(na1288_1), .IN1(~na172_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1975_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y62     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1289_1 ( .OUT(na1289_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na805_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1289_2 ( .OUT(na1289_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_10), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1289_6 ( .RAM_O1(na1289_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1289_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y61     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1290_4 ( .OUT(na1290_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na802_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1290_5 ( .OUT(na1290_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_11), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1290_6 ( .RAM_O2(na1290_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1290_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y61     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1291_1 ( .OUT(na1291_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na513_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1291_2 ( .OUT(na1291_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_12), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1291_6 ( .RAM_O1(na1291_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1291_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x88y76     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1292_1 ( .OUT(na1292_1), .IN1(~na177_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1976_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y60     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1293_4 ( .OUT(na1293_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na796_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1293_5 ( .OUT(na1293_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_13), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1293_6 ( .RAM_O2(na1293_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1293_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y60     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1294_1 ( .OUT(na1294_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na792_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1294_2 ( .OUT(na1294_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_14), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1294_6 ( .RAM_O1(na1294_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1294_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y59     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1295_4 ( .OUT(na1295_2_i), .IN1(na850_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1295_5 ( .OUT(na1295_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_15), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1295_6 ( .RAM_O2(na1295_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1295_2_i), .COMP_OUT(1'b0) );
// C_ORAND////      x90y79     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1296_1 ( .OUT(na1296_1), .IN1(~na182_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1977_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y59     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1297_1 ( .OUT(na1297_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na440_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1297_2 ( .OUT(na1297_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_16), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1297_6 ( .RAM_O1(na1297_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1297_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y58     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1298_4 ( .OUT(na1298_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na847_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1298_5 ( .OUT(na1298_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_17), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1298_6 ( .RAM_O2(na1298_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1298_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y58     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1299_1 ( .OUT(na1299_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na787_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1299_2 ( .OUT(na1299_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_18), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1299_6 ( .RAM_O1(na1299_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1299_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x90y78     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1300_1 ( .OUT(na1300_1), .IN1(~na187_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1978_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y57     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1301_4 ( .OUT(na1301_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na351_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1301_5 ( .OUT(na1301_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_19), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1301_6 ( .RAM_O2(na1301_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1301_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y57     80'h05_0018_00_0000_0C88_F5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1302_1 ( .OUT(na1302_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na270_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1302_2 ( .OUT(na1302_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_20), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1302_6 ( .RAM_O1(na1302_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1302_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y62     80'h0A_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1303_4 ( .OUT(na1303_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na727_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1303_5 ( .OUT(na1303_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_89), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1303_6 ( .RAM_O2(na1303_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1303_2_i), .COMP_OUT(1'b0) );
// C_ORAND////      x82y81     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1304_1 ( .OUT(na1304_1), .IN1(~na192_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1979_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x66y62     80'h05_0018_00_0000_0C88_F3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1305_1 ( .OUT(na1305_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na718_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1305_2 ( .OUT(na1305_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_90), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1305_6 ( .RAM_O1(na1305_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1305_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y61     80'h0A_0060_00_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1306_4 ( .OUT(na1306_2_i), .IN1(~na711_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1306_5 ( .OUT(na1306_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_91), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1306_6 ( .RAM_O2(na1306_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1306_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y61     80'h05_0018_00_0000_0C88_F5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1307_1 ( .OUT(na1307_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na702_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1307_2 ( .OUT(na1307_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_92), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1307_6 ( .RAM_O1(na1307_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1307_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x86y83     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1308_1 ( .OUT(na1308_1), .IN1(~na197_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1980_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x66y60     80'h0A_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1309_4 ( .OUT(na1309_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na693_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1309_5 ( .OUT(na1309_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_93), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1309_6 ( .RAM_O2(na1309_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1309_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y60     80'h05_0018_00_0000_0C88_F3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1310_1 ( .OUT(na1310_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na683_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1310_2 ( .OUT(na1310_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_94), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1310_6 ( .RAM_O1(na1310_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1310_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y59     80'h0A_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1311_4 ( .OUT(na1311_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na677_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1311_5 ( .OUT(na1311_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_95), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1311_6 ( .RAM_O2(na1311_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1311_2_i), .COMP_OUT(1'b0) );
// C_ORAND////      x92y79     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1312_1 ( .OUT(na1312_1), .IN1(~na202_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1983_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x66y59     80'h05_0018_00_0000_0C88_3FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1313_1 ( .OUT(na1313_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na671_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1313_2 ( .OUT(na1313_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_96), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1313_6 ( .RAM_O1(na1313_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1313_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y58     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1314_4 ( .OUT(na1314_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na838_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1314_5 ( .OUT(na1314_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_97), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1314_6 ( .RAM_O2(na1314_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1314_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y58     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1315_1 ( .OUT(na1315_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na655_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1315_2 ( .OUT(na1315_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_98), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1315_6 ( .RAM_O1(na1315_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1315_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x94y80     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1316_1 ( .OUT(na1316_1), .IN1(~na207_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1984_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x66y57     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1317_4 ( .OUT(na1317_2_i), .IN1(na833_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1317_5 ( .OUT(na1317_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_99), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1317_6 ( .RAM_O2(na1317_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1317_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y57     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1318_1 ( .OUT(na1318_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na641_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1318_2 ( .OUT(na1318_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1213_100), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1318_6 ( .RAM_O1(na1318_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1318_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x67y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1319_4 ( .OUT(na1319_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1319_6 ( .RAM_O2(na1319_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1319_2), .COMP_OUT(1'b0) );
// C_ORAND////      x92y80     80'h00_0018_00_0000_0888_3E57
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1320_1 ( .OUT(na1320_1), .IN1(~na212_1), .IN2(~na1228_2), .IN3(~na42_1), .IN4(1'b0), .IN5(na1985_2), .IN6(na1228_2), .IN7(1'b0),
                      .IN8(~na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x67y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1321_1 ( .OUT(na1321_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1321_6 ( .RAM_O1(na1321_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1321_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x67y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1322_4 ( .OUT(na1322_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1322_6 ( .RAM_O2(na1322_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1322_2), .COMP_OUT(1'b0) );
// C_AND////      x67y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1323_1 ( .OUT(na1323_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1323_6 ( .RAM_O1(na1323_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1323_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x65y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1324_4 ( .OUT(na1324_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1324_6 ( .RAM_O2(na1324_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1324_2), .COMP_OUT(1'b0) );
// C_AND////      x65y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1325_1 ( .OUT(na1325_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1325_6 ( .RAM_O1(na1325_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1325_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x84y53     80'h00_0018_00_0000_0888_1532
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1326_1 ( .OUT(na1326_1), .IN1(na1732_1), .IN2(~na1327_1), .IN3(1'b1), .IN4(~na348_2), .IN5(~na334_1), .IN6(1'b1), .IN7(~na336_1),
                      .IN8(~na348_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y66     80'h00_0018_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1327_1 ( .OUT(na1327_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na777_1), .IN6(na1932_2), .IN7(1'b0), .IN8(na102_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x65y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1328_4 ( .OUT(na1328_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1328_6 ( .RAM_O2(na1328_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1328_2), .COMP_OUT(1'b0) );
// C_ORAND////      x88y79     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1329_1 ( .OUT(na1329_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na314_2), .IN6(1'b0), .IN7(~na10_1), .IN8(na516_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x65y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1330_1 ( .OUT(na1330_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1330_6 ( .RAM_O1(na1330_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1330_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x82y77     80'h00_0018_00_0000_0C88_37FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1331_1 ( .OUT(na1331_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2073_2), .IN6(~na8_1), .IN7(1'b0), .IN8(~na1936_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y75     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1332_1 ( .OUT(na1332_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na316_1), .IN8(~na319_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x77y70     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1333_1 ( .OUT(na1333_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1937_2), .IN6(1'b0), .IN7(na406_1), .IN8(~na7_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x67y66     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1334_1 ( .OUT(na1334_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na240_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1334_6 ( .RAM_O1(na1334_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1334_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x59y65     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1335_4 ( .OUT(na1335_2), .IN1(1'b1), .IN2(na39_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1335_6 ( .RAM_O2(na1335_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1335_2), .COMP_OUT(1'b0) );
// C_MX2b////      x71y58     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1336_1 ( .OUT(na1336_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na952_1), .IN7(1'b0), .IN8(na984_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x76y47     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1337_1 ( .OUT(na1337_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na85_1), .IN6(1'b1), .IN7(~na83_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1338_4 ( .OUT(na1338_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1338_6 ( .RAM_O2(na1338_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1338_2), .COMP_OUT(1'b0) );
// C_AND////      x60y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1339_1 ( .OUT(na1339_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1339_6 ( .RAM_O1(na1339_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1339_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1340_4 ( .OUT(na1340_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1340_6 ( .RAM_O2(na1340_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1340_2), .COMP_OUT(1'b0) );
// C_AND///AND/      x93y49     80'h00_0078_00_0000_0C88_1FC3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1341_1 ( .OUT(na1341_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na346_1), .IN8(~na49_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1341_4 ( .OUT(na1341_2), .IN1(1'b1), .IN2(~na2021_2), .IN3(1'b1), .IN4(na44_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x81y52     80'h00_0018_00_0000_0888_F7D3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1342_1 ( .OUT(na1342_1), .IN1(1'b0), .IN2(~na342_1), .IN3(~na510_2), .IN4(na344_1), .IN5(~na1064_1), .IN6(~na1142_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1343_1 ( .OUT(na1343_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1343_6 ( .RAM_O1(na1343_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1343_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y70     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1344_4 ( .OUT(na1344_2), .IN1(na1062_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1344_6 ( .RAM_O2(na1344_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1344_2), .COMP_OUT(1'b0) );
// C_AND////      x60y70     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1345_1 ( .OUT(na1345_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1061_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1345_6 ( .RAM_O1(na1345_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1345_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x75y60     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1346_4 ( .OUT(na1346_2), .IN1(~na1347_1), .IN2(1'b1), .IN3(1'b1), .IN4(na350_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x77y63     80'h00_0018_00_0000_0888_7B73
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1347_1 ( .OUT(na1347_1), .IN1(1'b0), .IN2(~na352_1), .IN3(~na1355_1), .IN4(~na102_1), .IN5(na380_1), .IN6(~na101_1), .IN7(~na783_1),
                      .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x82y80     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1348_1 ( .OUT(na1348_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1349_1), .IN6(~na8_1), .IN7(~na369_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y77     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1349_1 ( .OUT(na1349_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na368_1), .IN6(~na367_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x83y76     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1350_1 ( .OUT(na1350_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1351_1), .IN6(~na8_1), .IN7(~na376_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x75y79     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1351_1 ( .OUT(na1351_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na375_1), .IN8(~na374_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x80y69     80'h00_0018_00_0000_0C88_75FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1352_1 ( .OUT(na1352_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na378_1), .IN6(1'b0), .IN7(~na1353_1), .IN8(~na7_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y69     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1353_1 ( .OUT(na1353_1), .IN1(1'b1), .IN2(na4_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na328_1), .IN8(~na325_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y69     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1354_4 ( .OUT(na1354_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1060_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1354_6 ( .RAM_O2(na1354_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1354_2), .COMP_OUT(1'b0) );
// C_MX2b////      x74y49     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1355_1 ( .OUT(na1355_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na952_2), .IN7(1'b0), .IN8(na984_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x86y59     80'h00_0078_00_0000_0CEE_0D70
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1356_1 ( .OUT(na1356_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1341_2), .IN6(na386_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1356_4 ( .OUT(na1356_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na862_1), .IN4(~na350_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y57     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1357_4 ( .OUT(na1357_2), .IN1(1'b1), .IN2(na929_1), .IN3(na346_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y69     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1358_1 ( .OUT(na1358_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1059_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1358_6 ( .RAM_O1(na1358_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1358_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x82y56     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1359_1 ( .OUT(na1359_1), .IN1(1'b1), .IN2(na1982_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1173_1), .IN6(na1160_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y68     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1360_4 ( .OUT(na1360_2), .IN1(na1058_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1360_6 ( .RAM_O2(na1360_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1360_2), .COMP_OUT(1'b0) );
// C_///AND/      x86y70     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1361_4 ( .OUT(na1361_2), .IN1(1'b1), .IN2(1'b1), .IN3(na247_2), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y79     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1362_4 ( .OUT(na1362_2), .IN1(~na399_1), .IN2(~na391_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y68     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1363_1 ( .OUT(na1363_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1363_6 ( .RAM_O1(na1363_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1363_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x87y80     80'h00_0018_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1364_1 ( .OUT(na1364_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na10_1), .IN8(~na396_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y76     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1365_1 ( .OUT(na1365_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1873_2), .IN5(~na395_1), .IN6(1'b0), .IN7(~na393_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x92y77     80'h00_0018_00_0000_0C88_EDFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1366_1 ( .OUT(na1366_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1875_2), .IN6(na1962_2), .IN7(na10_1), .IN8(na1956_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y67     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1367_4 ( .OUT(na1367_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1367_6 ( .RAM_O2(na1367_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1367_2), .COMP_OUT(1'b0) );
// C_AND////      x60y67     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1368_1 ( .OUT(na1368_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1368_6 ( .RAM_O1(na1368_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1368_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y66     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1369_4 ( .OUT(na1369_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1369_6 ( .RAM_O2(na1369_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1369_2), .COMP_OUT(1'b0) );
// C_MX2b////      x74y77     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1370_1 ( .OUT(na1370_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na406_1), .IN8(~na319_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1371_1 ( .OUT(na1371_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1371_6 ( .RAM_O1(na1371_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1371_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x92y71     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1372_1 ( .OUT(na1372_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na408_1), .IN7(1'b1), .IN8(na11_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1373_4 ( .OUT(na1373_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1373_6 ( .RAM_O2(na1373_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1373_2), .COMP_OUT(1'b0) );
// C_MX2b////      x76y49     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1374_1 ( .OUT(na1374_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na974_1), .IN6(1'b0), .IN7(na1006_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x84y61     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1375_4 ( .OUT(na1375_2), .IN1(na940_1), .IN2(1'b1), .IN3(na346_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x91y49     80'h00_0078_00_0000_0CEE_A533
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1376_1 ( .OUT(na1376_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1341_2), .IN6(1'b0), .IN7(na1377_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1376_4 ( .OUT(na1376_2), .IN1(1'b0), .IN2(~na1023_1), .IN3(1'b0), .IN4(~na350_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x84y51     80'h00_0018_00_0000_0888_DF37
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1377_1 ( .OUT(na1377_1), .IN1(~na1064_1), .IN2(~na1154_1), .IN3(1'b0), .IN4(~na415_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na510_2),
                      .IN8(na417_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1378_1 ( .OUT(na1378_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1378_6 ( .RAM_O1(na1378_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1378_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x88y66     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1379_4 ( .OUT(na1379_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1903_2), .IN4(~na250_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1380_4 ( .OUT(na1380_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1380_6 ( .RAM_O2(na1380_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1380_2), .COMP_OUT(1'b0) );
// C_AND////      x69y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1381_1 ( .OUT(na1381_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1381_6 ( .RAM_O1(na1381_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1381_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x82y76     80'h00_0018_00_0000_0C88_73FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1382_1 ( .OUT(na1382_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na419_1), .IN7(~na10_1), .IN8(~na1383_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y74     80'h00_0018_00_0040_0AAA_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1383_1 ( .OUT(na1383_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1873_2), .IN5(1'b0), .IN6(~na424_1), .IN7(1'b0), .IN8(~na423_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y77     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1384_1 ( .OUT(na1384_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na499_1), .IN6(~na8_1), .IN7(1'b0), .IN8(~na427_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1385_4 ( .OUT(na1385_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1385_6 ( .RAM_O2(na1385_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1385_2), .COMP_OUT(1'b0) );
// C_ORAND////      x77y69     80'h00_0018_00_0000_0C88_B3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1386_1 ( .OUT(na1386_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na430_1), .IN7(na375_1), .IN8(~na7_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1387_1 ( .OUT(na1387_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1387_6 ( .RAM_O1(na1387_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1387_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y70     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1388_4 ( .OUT(na1388_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1153_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1388_6 ( .RAM_O2(na1388_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1388_2), .COMP_OUT(1'b0) );
// C_MX2b////      x78y51     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1389_1 ( .OUT(na1389_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na974_2), .IN6(1'b0), .IN7(na1006_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y54     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1390_1 ( .OUT(na1390_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na944_1), .IN7(na346_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x73y59     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1391_4 ( .OUT(na1391_2), .IN1(na1341_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na436_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y70     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1392_1 ( .OUT(na1392_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1152_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1392_6 ( .RAM_O1(na1392_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1392_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x84y56     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1393_1 ( .OUT(na1393_1), .IN1(1'b1), .IN2(na1982_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1145_1), .IN6(na1162_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x81y56     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1394_4 ( .OUT(na1394_2), .IN1(1'b0), .IN2(~na1943_2), .IN3(1'b0), .IN4(~na876_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y65     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1395_4 ( .OUT(na1395_2), .IN1(1'b1), .IN2(na918_1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y54     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1396_1 ( .OUT(na1396_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na441_1), .IN6(1'b1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x80y59     80'h00_0078_00_0000_0C88_C5C3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1397_1 ( .OUT(na1397_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na444_1), .IN6(1'b1), .IN7(1'b1), .IN8(na102_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1397_4 ( .OUT(na1397_2), .IN1(1'b1), .IN2(~na453_1), .IN3(1'b1), .IN4(na102_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y69     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1398_4 ( .OUT(na1398_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1151_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1398_6 ( .RAM_O2(na1398_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1398_2), .COMP_OUT(1'b0) );
// C_AND////      x88y63     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1399_1 ( .OUT(na1399_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na443_1), .IN8(na11_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x78y77     80'h00_0018_00_0000_0C88_73FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1400_1 ( .OUT(na1400_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na446_1), .IN7(~na10_1), .IN8(~na1401_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x78y76     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1401_1 ( .OUT(na1401_1), .IN1(1'b1), .IN2(na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na284_1), .IN6(~na276_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x79y75     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1402_1 ( .OUT(na1402_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1934_2), .IN6(~na8_1), .IN7(1'b0), .IN8(~na449_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y69     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1403_1 ( .OUT(na1403_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1150_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1403_6 ( .RAM_O1(na1403_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1403_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y68     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1404_4 ( .OUT(na1404_2), .IN1(1'b1), .IN2(na1149_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1404_6 ( .RAM_O2(na1404_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1404_2), .COMP_OUT(1'b0) );
// C_AND////      x69y68     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1405_1 ( .OUT(na1405_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1405_6 ( .RAM_O1(na1405_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1405_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y67     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1406_4 ( .OUT(na1406_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1406_6 ( .RAM_O2(na1406_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1406_2), .COMP_OUT(1'b0) );
// C_///AND/      x90y59     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1407_4 ( .OUT(na1407_2), .IN1(na945_1), .IN2(1'b1), .IN3(na346_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x79y57     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1408_4 ( .OUT(na1408_2), .IN1(na1341_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na456_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y67     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1409_1 ( .OUT(na1409_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1409_6 ( .RAM_O1(na1409_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1409_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x80y56     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1410_1 ( .OUT(na1410_1), .IN1(1'b1), .IN2(na1982_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1146_1), .IN6(na1163_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x86y58     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1411_4 ( .OUT(na1411_2), .IN1(1'b0), .IN2(~na1025_1), .IN3(1'b0), .IN4(~na350_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y61     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1412_1 ( .OUT(na1412_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na918_2), .IN7(1'b1), .IN8(na49_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x81y77     80'h00_0018_00_0000_0C88_73FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1413_1 ( .OUT(na1413_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na463_2), .IN7(~na10_1), .IN8(~na1414_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y76     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1414_1 ( .OUT(na1414_1), .IN1(1'b1), .IN2(~na8_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na462_1), .IN8(~na358_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x78y80     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1415_1 ( .OUT(na1415_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1946_2), .IN6(~na8_1), .IN7(1'b0), .IN8(~na1954_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y66     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1416_4 ( .OUT(na1416_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1416_6 ( .RAM_O2(na1416_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1416_2), .COMP_OUT(1'b0) );
// C_ORAND////      x77y75     80'h00_0018_00_0000_0C88_37FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1417_1 ( .OUT(na1417_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2083_2), .IN6(~na8_1), .IN7(1'b0), .IN8(~na1955_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y75     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1418_1 ( .OUT(na1418_1), .IN1(1'b1), .IN2(na1871_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na371_1), .IN8(~na1948_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y66     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1419_1 ( .OUT(na1419_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1419_6 ( .RAM_O1(na1419_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1419_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x76y53     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1420_1 ( .OUT(na1420_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na978_2), .IN7(1'b0), .IN8(na1011_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x83y58     80'h00_0078_00_0000_0CEE_0D70
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1421_1 ( .OUT(na1421_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1341_2), .IN6(na474_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1421_4 ( .OUT(na1421_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na878_1), .IN4(~na350_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y57     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1422_4 ( .OUT(na1422_2), .IN1(1'b1), .IN2(na946_1), .IN3(na346_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y65     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1423_4 ( .OUT(na1423_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1423_6 ( .RAM_O2(na1423_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1423_2), .COMP_OUT(1'b0) );
// C_MX2b////      x76y56     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1424_1 ( .OUT(na1424_1), .IN1(1'b1), .IN2(na1982_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1147_1), .IN6(na1164_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y65     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1425_1 ( .OUT(na1425_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1425_6 ( .RAM_O1(na1425_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1425_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x87y65     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1426_4 ( .OUT(na1426_2), .IN1(na922_1), .IN2(1'b1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x81y73     80'h00_0018_00_0000_0C88_75FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1427_1 ( .OUT(na1427_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na480_1), .IN6(1'b0), .IN7(~na10_1), .IN8(~na1428_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x82y74     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1428_1 ( .OUT(na1428_1), .IN1(1'b1), .IN2(~na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na395_1), .IN6(~na397_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x87y77     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1429_1 ( .OUT(na1429_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1951_2), .IN6(~na8_1), .IN7(~na484_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x62y72     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1430_4 ( .OUT(na1430_2_i), .IN1(na827_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1430_5 ( .OUT(na1430_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_21), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1430_6 ( .RAM_O2(na1430_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1430_2_i), .COMP_OUT(1'b0) );
// C_ORAND////      x91y71     80'h00_0018_00_0000_0C88_B3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1431_1 ( .OUT(na1431_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1952_2), .IN7(na486_1), .IN8(~na11_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y73     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1432_1 ( .OUT(na1432_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na486_1), .IN8(na11_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x62y72     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1433_1 ( .OUT(na1433_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na824_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1433_2 ( .OUT(na1433_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_22), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1433_6 ( .RAM_O1(na1433_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1433_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x72y53     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1434_1 ( .OUT(na1434_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na980_1), .IN6(1'b0), .IN7(na1013_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y50     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1435_1 ( .OUT(na1435_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(~na489_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x62y71     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1436_4 ( .OUT(na1436_2_i), .IN1(1'b1), .IN2(na616_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1436_5 ( .OUT(na1436_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_23), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1436_6 ( .RAM_O2(na1436_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1436_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x72y56     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1437_1 ( .OUT(na1437_1), .IN1(1'b1), .IN2(~na1982_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1166_1), .IN6(na1148_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x92y57     80'h00_0060_00_0000_0C0E_FF53
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1438_4 ( .OUT(na1438_2), .IN1(1'b0), .IN2(~na946_2), .IN3(~na346_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y57     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1439_4 ( .OUT(na1439_2), .IN1(1'b1), .IN2(na1943_2), .IN3(1'b1), .IN4(na1027_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x91y65     80'h00_0018_00_0000_0C88_B3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1440_1 ( .OUT(na1440_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1952_2), .IN7(na495_1), .IN8(~na11_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y67     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1441_1 ( .OUT(na1441_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na495_1), .IN8(na11_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x62y71     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1442_1 ( .OUT(na1442_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na821_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1442_2 ( .OUT(na1442_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_24), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1442_6 ( .RAM_O1(na1442_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1442_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x84y78     80'h00_0018_00_0000_0C88_75FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1443_1 ( .OUT(na1443_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na498_1), .IN6(1'b0), .IN7(~na10_1), .IN8(~na1444_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y74     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1444_1 ( .OUT(na1444_1), .IN1(1'b1), .IN2(na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na420_1), .IN6(~na424_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y78     80'h00_0018_00_0000_0C88_37FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1445_1 ( .OUT(na1445_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1446_1), .IN6(~na8_1), .IN7(1'b0), .IN8(~na503_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x69y77     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1446_1 ( .OUT(na1446_1), .IN1(1'b1), .IN2(~na1871_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na371_1), .IN8(~na374_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y72     80'h0A_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1447_4 ( .OUT(na1447_2_i), .IN1(1'b1), .IN2(na594_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1447_5 ( .OUT(na1447_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_25), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1447_6 ( .RAM_O2(na1447_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1447_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x70y51     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1448_1 ( .OUT(na1448_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na980_2), .IN6(1'b0), .IN7(na1013_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x86y58     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1449_1 ( .OUT(na1449_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na948_1), .IN6(1'b1), .IN7(na346_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x97y48     80'h00_0078_00_0000_0CEE_0D33
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1450_1 ( .OUT(na1450_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1341_2), .IN6(na1451_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1450_4 ( .OUT(na1450_2), .IN1(1'b0), .IN2(~na1943_2), .IN3(1'b0), .IN4(~na880_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x87y48     80'h00_0018_00_0000_0888_DFDC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1451_1 ( .OUT(na1451_1), .IN1(1'b0), .IN2(na512_1), .IN3(~na510_1), .IN4(na1959_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na510_2),
                      .IN8(na511_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y72     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1452_1 ( .OUT(na1452_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na581_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1452_2 ( .OUT(na1452_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_26), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1452_6 ( .RAM_O1(na1452_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1452_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x85y65     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1453_4 ( .OUT(na1453_2), .IN1(1'b1), .IN2(na924_1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y71     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1454_4 ( .OUT(na1454_2_i), .IN1(na568_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1454_5 ( .OUT(na1454_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_27), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1454_6 ( .RAM_O2(na1454_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1454_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y71     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1455_1 ( .OUT(na1455_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na812_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1455_2 ( .OUT(na1455_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_28), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1455_6 ( .RAM_O1(na1455_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1455_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x71y59     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1456_4 ( .OUT(na1456_2), .IN1(1'b1), .IN2(~na509_1), .IN3(na2029_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y56     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1457_4 ( .OUT(na1457_2), .IN1(na1942_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1458_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y66     80'h00_0018_00_0000_0888_7BB3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1458_1 ( .OUT(na1458_1), .IN1(1'b0), .IN2(~na514_1), .IN3(na518_1), .IN4(~na102_1), .IN5(na517_1), .IN6(~na101_1), .IN7(~na797_1),
                      .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y70     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1459_4 ( .OUT(na1459_2_i), .IN1(na809_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1459_5 ( .OUT(na1459_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_29), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1459_6 ( .RAM_O2(na1459_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1459_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x82y73     80'h00_0018_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1460_1 ( .OUT(na1460_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na10_1), .IN4(1'b1), .IN5(1'b0), .IN6(na283_1), .IN7(1'b0), .IN8(na516_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y54     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1461_1 ( .OUT(na1461_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na948_2), .IN6(1'b1), .IN7(na346_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x90y49     80'h00_0018_00_0000_0C88_BAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1462_1 ( .OUT(na1462_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b0), .IN7(na521_1), .IN8(~na523_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y70     80'h05_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1463_1 ( .OUT(na1463_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na805_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1463_2 ( .OUT(na1463_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_30), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1463_6 ( .RAM_O1(na1463_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1463_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x87y57     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1464_1 ( .OUT(na1464_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1029_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na350_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y62     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1465_4 ( .OUT(na1465_2), .IN1(1'b1), .IN2(na924_2), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y55     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1466_4 ( .OUT(na1466_2), .IN1(1'b1), .IN2(na1063_1), .IN3(1'b1), .IN4(~na344_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x89y79     80'h00_0018_00_0000_0C88_E7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1467_1 ( .OUT(na1467_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1875_2), .IN6(~na1469_1), .IN7(na10_1),
                      .IN8(na1348_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y69     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1468_4 ( .OUT(na1468_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na802_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1468_5 ( .OUT(na1468_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_31), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1468_6 ( .RAM_O2(na1468_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1468_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x79y82     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1469_1 ( .OUT(na1469_1), .IN1(1'b1), .IN2(na8_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na361_1), .IN8(~na358_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x91y68     80'h00_0018_00_0000_0C88_B3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1470_1 ( .OUT(na1470_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1952_2), .IN7(na482_1), .IN8(~na11_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y73     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1471_1 ( .OUT(na1471_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na482_1), .IN8(na11_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y53     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1472_1 ( .OUT(na1472_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na982_2), .IN7(1'b0), .IN8(na1015_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y52     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1473_4 ( .OUT(na1473_2), .IN1(na1341_2), .IN2(1'b1), .IN3(~na531_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y69     80'h05_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1474_1 ( .OUT(na1474_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na513_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1474_2 ( .OUT(na1474_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_32), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1474_6 ( .RAM_O1(na1474_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1474_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y68     80'h0A_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1475_4 ( .OUT(na1475_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na796_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1475_5 ( .OUT(na1475_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_33), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1475_6 ( .RAM_O2(na1475_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1475_2_i), .COMP_OUT(1'b0) );
// C_OR////      x88y57     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1476_1 ( .OUT(na1476_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na882_1), .IN8(~na350_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y59     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1477_1 ( .OUT(na1477_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na926_1), .IN6(1'b1), .IN7(1'b1), .IN8(na49_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y68     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1478_1 ( .OUT(na1478_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na792_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1478_2 ( .OUT(na1478_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_34), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1478_6 ( .RAM_O1(na1478_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1478_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x86y79     80'h00_0018_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1479_1 ( .OUT(na1479_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na10_1), .IN4(1'b1), .IN5(1'b0), .IN6(na1950_2), .IN7(1'b0), .IN8(na538_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y67     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1480_4 ( .OUT(na1480_2_i), .IN1(na850_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1480_5 ( .OUT(na1480_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_35), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1480_6 ( .RAM_O2(na1480_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1480_2_i), .COMP_OUT(1'b0) );
// C_AND////      x87y65     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1481_1 ( .OUT(na1481_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na466_1), .IN8(na11_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y61     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1482_1 ( .OUT(na1482_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na953_1), .IN6(1'b0), .IN7(na985_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x89y49     80'h00_0018_00_0000_0C88_BAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1483_1 ( .OUT(na1483_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b0), .IN7(na521_1), .IN8(~na544_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y67     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1484_1 ( .OUT(na1484_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na440_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1484_2 ( .OUT(na1484_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_36), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1484_6 ( .RAM_O1(na1484_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1484_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x97y56     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1485_1 ( .OUT(na1485_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na950_2), .IN7(na346_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x98y53     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1486_1 ( .OUT(na1486_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1031_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na350_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y67     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1487_4 ( .OUT(na1487_2), .IN1(na926_2), .IN2(1'b1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x79y49     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1488_1 ( .OUT(na1488_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1063_1), .IN7(1'b1), .IN8(~na417_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y73     80'h00_0018_00_0000_0888_CF7E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1489_1 ( .OUT(na1489_1), .IN1(na1384_1), .IN2(na1876_2), .IN3(~na10_1), .IN4(~na1490_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                      .IN8(na11_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y78     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1490_1 ( .OUT(na1490_1), .IN1(1'b1), .IN2(~na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na420_1), .IN6(~na421_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x64y66     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1491_4 ( .OUT(na1491_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na847_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1491_5 ( .OUT(na1491_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_37), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1491_6 ( .RAM_O2(na1491_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1491_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x64y66     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1492_1 ( .OUT(na1492_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na787_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1492_2 ( .OUT(na1492_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_38), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1492_6 ( .RAM_O1(na1492_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1492_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x64y65     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1493_4 ( .OUT(na1493_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na351_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1493_5 ( .OUT(na1493_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_39), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1493_6 ( .RAM_O2(na1493_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1493_2_i), .COMP_OUT(1'b0) );
// C_AND////      x85y65     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1494_1 ( .OUT(na1494_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1877_2), .IN7(1'b1), .IN8(~na447_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y53     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1495_1 ( .OUT(na1495_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na953_2), .IN6(1'b0), .IN7(na985_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x64y65     80'h05_0018_00_0000_0C88_F5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1496_1 ( .OUT(na1496_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na270_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1496_2 ( .OUT(na1496_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_40), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1496_6 ( .RAM_O1(na1496_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1496_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y70     80'h0A_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1497_4 ( .OUT(na1497_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na727_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1497_5 ( .OUT(na1497_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_109), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1497_6 ( .RAM_O2(na1497_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1497_2_i), .COMP_OUT(1'b0) );
// C_AND////      x98y55     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1498_1 ( .OUT(na1498_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na930_1), .IN6(1'b1), .IN7(na346_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x89y53     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1499_1 ( .OUT(na1499_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1943_2), .IN7(1'b0), .IN8(~na853_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y62     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1500_4 ( .OUT(na1500_2), .IN1(1'b1), .IN2(na928_1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y75     80'h00_0018_00_0000_0888_CF7E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1501_1 ( .OUT(na1501_1), .IN1(na1402_1), .IN2(na1876_2), .IN3(~na10_1), .IN4(~na1502_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                      .IN8(na11_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y80     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1502_1 ( .OUT(na1502_1), .IN1(1'b1), .IN2(~na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na291_1), .IN6(~na300_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x66y70     80'h05_0018_00_0000_0C88_F3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1503_1 ( .OUT(na1503_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na718_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1503_2 ( .OUT(na1503_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_110), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1503_6 ( .RAM_O1(na1503_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1503_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y69     80'h0A_0060_00_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1504_4 ( .OUT(na1504_2_i), .IN1(~na711_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1504_5 ( .OUT(na1504_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_111), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1504_6 ( .RAM_O2(na1504_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1504_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x77y60     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1505_1 ( .OUT(na1505_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na955_1), .IN7(1'b0), .IN8(na987_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y59     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1506_4 ( .OUT(na1506_2), .IN1(1'b1), .IN2(na567_1), .IN3(na2029_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x89y52     80'h00_0018_00_0000_0CEE_A500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1507_1 ( .OUT(na1507_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1341_2), .IN6(1'b0), .IN7(na564_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y58     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1508_1 ( .OUT(na1508_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na931_1), .IN7(na346_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x66y69     80'h05_0018_00_0000_0C88_F5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1509_1 ( .OUT(na1509_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na702_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1509_2 ( .OUT(na1509_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_112), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1509_6 ( .RAM_O1(na1509_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1509_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y68     80'h0A_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1510_4 ( .OUT(na1510_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na693_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1510_5 ( .OUT(na1510_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_113), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1510_6 ( .RAM_O2(na1510_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1510_2_i), .COMP_OUT(1'b0) );
// C_OR////      x93y53     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1511_1 ( .OUT(na1511_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1033_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na350_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y71     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1512_4 ( .OUT(na1512_2), .IN1(1'b1), .IN2(na928_2), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y54     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1513_1 ( .OUT(na1513_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na569_1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x66y68     80'h05_0018_00_0000_0C88_F3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1514_1 ( .OUT(na1514_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na683_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1514_2 ( .OUT(na1514_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_114), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1514_6 ( .RAM_O1(na1514_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1514_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x83y71     80'h00_0018_00_0000_0888_CFD3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1515_1 ( .OUT(na1515_1), .IN1(1'b0), .IN2(~na571_2), .IN3(~na10_1), .IN4(na1415_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0), .IN8(na11_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/RAM_I2      x66y67     80'h0A_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1516_4 ( .OUT(na1516_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na677_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1516_5 ( .OUT(na1516_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_115), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1516_6 ( .RAM_O2(na1516_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1516_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y67     80'h05_0018_00_0000_0C88_3FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1517_1 ( .OUT(na1517_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na671_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1517_2 ( .OUT(na1517_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_116), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1517_6 ( .RAM_O1(na1517_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1517_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y66     80'h0A_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1518_4 ( .OUT(na1518_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na838_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1518_5 ( .OUT(na1518_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_117), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1518_6 ( .RAM_O2(na1518_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1518_2_i), .COMP_OUT(1'b0) );
// C_AND/RAM_I1///      x66y66     80'h05_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1519_1 ( .OUT(na1519_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na655_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1519_2 ( .OUT(na1519_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_118), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1519_6 ( .RAM_O1(na1519_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1519_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/RAM_I2      x66y65     80'h0A_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1520_4 ( .OUT(na1520_2_i), .IN1(na833_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1520_5 ( .OUT(na1520_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_119), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1520_6 ( .RAM_O2(na1520_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1520_2_i), .COMP_OUT(1'b0) );
// C_MX2b////      x74y55     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1521_1 ( .OUT(na1521_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na955_2), .IN7(1'b0), .IN8(na987_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y57     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1522_4 ( .OUT(na1522_2), .IN1(1'b1), .IN2(1'b1), .IN3(na855_1), .IN4(na350_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x95y52     80'h00_0060_00_0000_0C0E_FF0D
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1523_4 ( .OUT(na1523_2), .IN1(~na1341_2), .IN2(na578_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y59     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1524_1 ( .OUT(na1524_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na932_1), .IN6(1'b1), .IN7(na346_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/RAM_I1///      x66y65     80'h05_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1525_1 ( .OUT(na1525_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na641_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0011)) 
           _a1525_2 ( .OUT(na1525_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na1214_120), .CP_O(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1525_6 ( .RAM_O1(na1525_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1525_1_i),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x67y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1526_4 ( .OUT(na1526_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1526_6 ( .RAM_O2(na1526_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1526_2), .COMP_OUT(1'b0) );
// C_///OR/      x90y55     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1527_4 ( .OUT(na1527_2), .IN1(~na1064_1), .IN2(~na567_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x82y72     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1528_4 ( .OUT(na1528_2), .IN1(na909_1), .IN2(1'b1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y62     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1529_1 ( .OUT(na1529_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na582_1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x67y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1530_1 ( .OUT(na1530_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1530_6 ( .RAM_O1(na1530_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1530_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x87y75     80'h00_0018_00_0000_0888_CF7E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1531_1 ( .OUT(na1531_1), .IN1(na1429_1), .IN2(na1876_2), .IN3(~na10_1), .IN4(~na1532_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                      .IN8(na11_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x80y82     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1532_1 ( .OUT(na1532_1), .IN1(1'b1), .IN2(~na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na398_1), .IN6(~na401_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x67y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1533_4 ( .OUT(na1533_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1533_6 ( .RAM_O2(na1533_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1533_2), .COMP_OUT(1'b0) );
// C_AND////      x67y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1534_1 ( .OUT(na1534_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1534_6 ( .RAM_O1(na1534_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1534_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x65y72     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1535_4 ( .OUT(na1535_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1535_6 ( .RAM_O2(na1535_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1535_2), .COMP_OUT(1'b0) );
// C_ORAND////      x90y81     80'h00_0018_00_0000_0C88_DEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1536_1 ( .OUT(na1536_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1875_2), .IN6(na1350_1), .IN7(~na10_1), .IN8(na1348_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y59     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1537_1 ( .OUT(na1537_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na957_1), .IN6(1'b0), .IN7(na989_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y51     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1538_1 ( .OUT(na1538_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na590_1), .IN6(na2076_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x65y72     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1539_1 ( .OUT(na1539_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1539_6 ( .RAM_O1(na1539_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1539_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x65y71     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1540_4 ( .OUT(na1540_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1540_6 ( .RAM_O2(na1540_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1540_2), .COMP_OUT(1'b0) );
// C_OR////      x89y62     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1541_1 ( .OUT(na1541_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na567_1), .IN7(1'b0), .IN8(~na1065_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y71     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1542_4 ( .OUT(na1542_2), .IN1(na909_2), .IN2(1'b1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x97y60     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1543_1 ( .OUT(na1543_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na933_1), .IN7(~na346_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y53     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1544_1 ( .OUT(na1544_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1035_1), .IN7(1'b1), .IN8(na350_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y58     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1545_1 ( .OUT(na1545_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na595_1), .IN6(1'b1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x65y71     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1546_1 ( .OUT(na1546_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1546_6 ( .RAM_O1(na1546_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1546_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x87y73     80'h00_0018_00_0000_0888_CFE7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1547_1 ( .OUT(na1547_1), .IN1(~na1875_2), .IN2(~na1548_1), .IN3(na10_1), .IN4(na1445_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                      .IN8(na11_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x79y78     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1548_1 ( .OUT(na1548_1), .IN1(1'b1), .IN2(na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na499_1), .IN6(~na421_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y59     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1553_1 ( .OUT(na1553_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na957_2), .IN6(1'b0), .IN7(na989_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x67y57     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1555_4 ( .OUT(na1555_2), .IN1(1'b1), .IN2(na1063_1), .IN3(1'b1), .IN4(~na511_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x91y60     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1556_4 ( .OUT(na1556_2), .IN1(1'b0), .IN2(~na1943_2), .IN3(1'b0), .IN4(~na857_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y57     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1557_1 ( .OUT(na1557_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na911_1), .IN7(1'b1), .IN8(na49_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x95y73     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1558_4 ( .OUT(na1558_2), .IN1(~na934_1), .IN2(1'b0), .IN3(~na346_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x98y55     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1559_4 ( .OUT(na1559_2), .IN1(1'b1), .IN2(na567_1), .IN3(1'b1), .IN4(na1066_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y57     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1561_1 ( .OUT(na1561_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na959_1), .IN7(1'b0), .IN8(na991_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y50     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1563_4 ( .OUT(na1563_2), .IN1(na1064_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1150_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x95y55     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1564_1 ( .OUT(na1564_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1037_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na350_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y71     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1565_4 ( .OUT(na1565_2), .IN1(1'b1), .IN2(na911_2), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x91y66     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1566_1 ( .OUT(na1566_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na935_1), .IN7(~na346_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y58     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1567_1 ( .OUT(na1567_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na567_1), .IN7(1'b1), .IN8(na1067_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x97y58     80'h00_0078_00_0000_0C88_C3AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1568_1 ( .OUT(na1568_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1569_1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1568_4 ( .OUT(na1568_2), .IN1(na936_1), .IN2(1'b1), .IN3(na346_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x81y62     80'h00_0018_00_0000_0888_3F14
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1569_1 ( .OUT(na1569_1), .IN1(~na1570_1), .IN2(na1574_2), .IN3(~na620_1), .IN4(~na617_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na617_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x85y71     80'h00_0018_00_0000_0C88_34FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1570_1 ( .OUT(na1570_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1531_1), .IN6(na101_1), .IN7(1'b1), .IN8(~na586_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x67y66     80'h00_0060_00_0000_0C0E_FFD5
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1574_4 ( .OUT(na1574_2), .IN1(~na84_1), .IN2(1'b0), .IN3(~na1436_2), .IN4(na24_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y63     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1576_1 ( .OUT(na1576_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na959_2), .IN7(1'b0), .IN8(na991_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y51     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1577_1 ( .OUT(na1577_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na859_1), .IN8(na350_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x86y52     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1580_4 ( .OUT(na1580_2), .IN1(na1064_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1151_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x91y57     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1581_1 ( .OUT(na1581_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na567_1), .IN7(1'b0), .IN8(~na1068_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y68     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1582_4 ( .OUT(na1582_2), .IN1(na913_1), .IN2(1'b1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x84y69     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1584_1 ( .OUT(na1584_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na961_1), .IN6(1'b0), .IN7(na993_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x84y63     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1585_4 ( .OUT(na1585_2), .IN1(1'b1), .IN2(na937_1), .IN3(na346_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y52     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1588_4 ( .OUT(na1588_2), .IN1(na1064_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1152_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x94y55     80'h00_0018_00_0000_0CEE_7000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1589_1 ( .OUT(na1589_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1039_1), .IN8(~na350_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x77y64     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1590_4 ( .OUT(na1590_2), .IN1(1'b1), .IN2(na567_1), .IN3(1'b1), .IN4(na1069_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x73y65     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1592_1 ( .OUT(na1592_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na961_2), .IN6(1'b0), .IN7(na993_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y54     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1593_1 ( .OUT(na1593_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1943_2), .IN7(1'b1), .IN8(na861_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y52     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1596_4 ( .OUT(na1596_2), .IN1(na1064_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1153_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x91y64     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1597_1 ( .OUT(na1597_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na938_1), .IN6(1'b0), .IN7(~na346_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y67     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1598_4 ( .OUT(na1598_2), .IN1(1'b1), .IN2(na915_1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x92y65     80'h00_0078_00_0000_0C88_CCAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1599_1 ( .OUT(na1599_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na915_2), .IN7(1'b1), .IN8(na49_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1599_4 ( .OUT(na1599_2), .IN1(1'b1), .IN2(na939_1), .IN3(na346_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y67     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1603_1 ( .OUT(na1603_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na964_1), .IN7(1'b0), .IN8(na996_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y50     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1606_4 ( .OUT(na1606_2), .IN1(na1064_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1155_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x95y54     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1607_1 ( .OUT(na1607_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1041_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na350_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y57     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1608_1 ( .OUT(na1608_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1058_2), .IN6(na567_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y67     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1612_1 ( .OUT(na1612_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na964_2), .IN7(1'b0), .IN8(na996_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y50     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1614_4 ( .OUT(na1614_2), .IN1(na1156_1), .IN2(1'b1), .IN3(na2031_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x89y58     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1615_4 ( .OUT(na1615_2), .IN1(~na1059_2), .IN2(~na567_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y61     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1616_1 ( .OUT(na1616_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na917_1), .IN6(1'b1), .IN7(1'b1), .IN8(na49_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x94y66     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1617_1 ( .OUT(na1617_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na941_1), .IN6(1'b0), .IN7(~na346_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x99y51     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1618_1 ( .OUT(na1618_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na864_1), .IN8(na350_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x90y57     80'h00_0078_00_0000_0C88_4FAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1619_1 ( .OUT(na1619_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na656_1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1619_4 ( .OUT(na1619_2), .IN1(1'b1), .IN2(na567_1), .IN3(na1060_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x74y65     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1623_1 ( .OUT(na1623_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na966_1), .IN6(1'b0), .IN7(na998_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y56     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1624_1 ( .OUT(na1624_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1943_2), .IN7(1'b1), .IN8(na1043_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y54     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1626_4 ( .OUT(na1626_2), .IN1(na1064_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1157_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x87y77     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1630_4 ( .OUT(na1630_2), .IN1(1'b1), .IN2(~na500_1), .IN3(1'b1), .IN4(na11_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y63     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1631_1 ( .OUT(na1631_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na966_2), .IN6(1'b0), .IN7(na998_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y58     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1632_4 ( .OUT(na1632_2), .IN1(na1061_2), .IN2(na567_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y52     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1635_1 ( .OUT(na1635_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1158_1), .IN6(1'b1), .IN7(na2031_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x88y60     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1636_4 ( .OUT(na1636_2), .IN1(1'b0), .IN2(~na1943_2), .IN3(1'b0), .IN4(~na866_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y63     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1637_1 ( .OUT(na1637_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na920_1), .IN7(1'b1), .IN8(na49_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x68y73     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1642_1 ( .OUT(na1642_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na968_1), .IN7(1'b0), .IN8(na1000_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x71y64     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1643_4 ( .OUT(na1643_2), .IN1(~na1064_1), .IN2(~na1159_1), .IN3(~na612_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x72y73     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1651_1 ( .OUT(na1651_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na968_2), .IN7(1'b0), .IN8(na1000_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x75y60     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1652_1 ( .OUT(na1652_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1064_1), .IN6(~na1160_1), .IN7(~na612_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x74y57     80'h00_0018_00_0000_0888_5515
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1657_1 ( .OUT(na1657_1), .IN1(~na689_1), .IN2(1'b1), .IN3(~na684_1), .IN4(~na687_1), .IN5(~na1658_2), .IN6(1'b1), .IN7(~na684_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x75y61     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1658_4 ( .OUT(na1658_2), .IN1(~na469_1), .IN2(1'b1), .IN3(1'b1), .IN4(na102_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x73y60     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1662_1 ( .OUT(na1662_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1064_1), .IN6(~na1161_1), .IN7(~na612_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x74y51     80'h00_0018_00_0000_0888_331A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1667_1 ( .OUT(na1667_1), .IN1(na1671_1), .IN2(1'b1), .IN3(~na695_1), .IN4(~na1668_1), .IN5(1'b1), .IN6(~na698_1), .IN7(1'b1),
                      .IN8(~na1668_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x80y66     80'h00_0078_00_0000_0C88_F4CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1668_1 ( .OUT(na1668_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na444_1), .IN6(na101_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1668_4 ( .OUT(na1668_2), .IN1(1'b1), .IN2(na1909_2), .IN3(1'b1), .IN4(na1673_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x71y59     80'h00_0018_00_0000_0CEE_7A00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1671_1 ( .OUT(na1671_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na34_1), .IN6(1'b0), .IN7(~na1905_2), .IN8(~na1510_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x76y64     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1673_1 ( .OUT(na1673_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na970_2), .IN6(1'b0), .IN7(na1002_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x91y54     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1676_4 ( .OUT(na1676_2), .IN1(~na1064_1), .IN2(~na1162_1), .IN3(~na612_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x84y59     80'h00_0018_00_0000_0EEE_0EEC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1681_1 ( .OUT(na1681_1), .IN1(1'b0), .IN2(na1682_2), .IN3(na706_1), .IN4(na708_1), .IN5(na1683_1), .IN6(na1682_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x81y70     80'h00_0078_00_0000_0C88_3C4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1682_1 ( .OUT(na1682_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na101_1), .IN7(1'b1), .IN8(~na418_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1682_4 ( .OUT(na1682_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na707_1), .IN4(na102_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x83y61     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1683_1 ( .OUT(na1683_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na431_1), .IN6(1'b1), .IN7(1'b1), .IN8(na102_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x89y54     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1687_4 ( .OUT(na1687_2), .IN1(~na1064_1), .IN2(~na1163_1), .IN3(~na612_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x76y65     80'h00_0018_00_0000_0888_775B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1692_1 ( .OUT(na1692_1), .IN1(na1362_2), .IN2(~na101_1), .IN3(~na714_1), .IN4(1'b0), .IN5(~na1695_1), .IN6(~na1909_2), .IN7(~na843_1),
                      .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y75     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1695_1 ( .OUT(na1695_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b0), .IN6(na972_2), .IN7(1'b0), .IN8(na1004_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x81y66     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1698_1 ( .OUT(na1698_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1064_1), .IN6(~na1164_1), .IN7(~na612_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x82y64     80'h00_0060_00_0000_0C0E_FFAB
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1703_4 ( .OUT(na1703_2), .IN1(na364_1), .IN2(~na101_1), .IN3(na782_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x84y71     80'h00_0078_00_0000_0C88_C5CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1705_1 ( .OUT(na1705_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na380_1), .IN6(1'b1), .IN7(1'b1), .IN8(na102_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1705_4 ( .OUT(na1705_2), .IN1(1'b1), .IN2(na1710_1), .IN3(1'b1), .IN4(na102_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x67y60     80'h00_0018_00_0000_0CEE_3D00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1708_1 ( .OUT(na1708_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na84_1), .IN6(na37_1), .IN7(1'b0), .IN8(~na1503_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x77y68     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1710_1 ( .OUT(na1710_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na975_1), .IN6(1'b0), .IN7(na1007_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y52     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1712_1 ( .OUT(na1712_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1064_1), .IN6(~na1166_1), .IN7(~na612_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x82y57     80'h00_0018_00_0000_0888_5435
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1715_1 ( .OUT(na1715_1), .IN1(~na732_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1717_1), .IN5(~na1718_1), .IN6(na731_1), .IN7(~na728_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y66     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1717_1 ( .OUT(na1717_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1911_2), .IN7(1'b1), .IN8(~na330_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x73y59     80'h00_0018_00_0000_0C88_DAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1718_1 ( .OUT(na1718_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na85_1), .IN6(1'b0), .IN7(~na1898_2), .IN8(na1497_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x69y79     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1720_1 ( .OUT(na1720_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na335_1), .IN5(na975_2), .IN6(1'b0), .IN7(na1007_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x77y70     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1721_4 ( .OUT(na1721_2), .IN1(~na1064_1), .IN2(~na1167_1), .IN3(~na612_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x83y74     80'h00_0018_00_0040_0AA2_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1730_1 ( .OUT(na1730_1), .IN1(1'b1), .IN2(1'b1), .IN3(na10_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na283_1), .IN7(1'b0), .IN8(na776_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x67y56     80'h00_0018_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1731_1 ( .OUT(na1731_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na4_1), .IN7(na1496_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x77y67     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1732_1 ( .OUT(na1732_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1064_1), .IN6(~na778_1), .IN7(~na2029_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x82y71     80'h00_0060_00_0000_0C08_FF73
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1734_4 ( .OUT(na1734_2), .IN1(1'b0), .IN2(~na357_1), .IN3(~na10_1), .IN4(~na781_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y73     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1735_4 ( .OUT(na1735_2), .IN1(1'b1), .IN2(1'b1), .IN3(na10_1), .IN4(na781_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y52     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1738_4 ( .OUT(na1738_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1739_1), .IN4(na350_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y53     80'h00_0018_00_0000_0888_7753
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1739_1 ( .OUT(na1739_1), .IN1(1'b0), .IN2(~na390_1), .IN3(~na407_2), .IN4(1'b0), .IN5(~na785_1), .IN6(~na2033_2), .IN7(~na1374_1),
                      .IN8(~na102_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y51     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1741_4 ( .OUT(na1741_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1742_1), .IN4(na350_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x88y55     80'h00_0018_00_0000_0888_7773
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1742_1 ( .OUT(na1742_1), .IN1(1'b0), .IN2(~na485_1), .IN3(~na479_1), .IN4(~na102_2), .IN5(~na790_1), .IN6(~na2033_2), .IN7(~na1434_1),
                      .IN8(~na102_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y55     80'h00_0018_00_0000_0C88_C8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1743_1 ( .OUT(na1743_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1941_2), .IN6(na2033_2), .IN7(1'b1), .IN8(na793_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y53     80'h00_0018_00_0000_0888_3C34
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1745_1 ( .OUT(na1745_1), .IN1(~na1453_2), .IN2(na1450_1), .IN3(1'b1), .IN4(~na1449_1), .IN5(1'b1), .IN6(na1450_2), .IN7(1'b1),
                      .IN8(~na350_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y56     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1750_1 ( .OUT(na1750_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1751_1), .IN6(1'b1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y57     80'h00_0018_00_0000_0888_77B5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1751_1 ( .OUT(na1751_1), .IN1(~na528_2), .IN2(1'b0), .IN3(na525_1), .IN4(~na102_2), .IN5(~na800_1), .IN6(~na2033_2), .IN7(~na1472_1),
                      .IN8(~na102_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y53     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1753_4 ( .OUT(na1753_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1754_1), .IN4(na350_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y55     80'h00_0018_00_0000_0888_7755
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1754_1 ( .OUT(na1754_1), .IN1(~na539_1), .IN2(1'b0), .IN3(~na535_1), .IN4(1'b0), .IN5(~na2032_2), .IN6(~na803_1), .IN7(~na1482_1),
                      .IN8(~na102_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y50     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1756_1 ( .OUT(na1756_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1341_2), .IN6(1'b1), .IN7(~na551_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x87y51     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1757_1 ( .OUT(na1757_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1758_1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x83y56     80'h00_0018_00_0000_0888_7753
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1758_1 ( .OUT(na1758_1), .IN1(1'b0), .IN2(~na545_2), .IN3(~na549_1), .IN4(1'b0), .IN5(~na806_1), .IN6(~na2033_2), .IN7(~na1495_1),
                      .IN8(~na102_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y59     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1760_1 ( .OUT(na1760_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1761_1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x81y64     80'h00_0018_00_0000_0888_775B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1761_1 ( .OUT(na1761_1), .IN1(na1963_2), .IN2(~na101_1), .IN3(~na557_2), .IN4(1'b0), .IN5(~na1908_2), .IN6(~na1505_1), .IN7(~na810_1),
                      .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y56     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1766_4 ( .OUT(na1766_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1767_1), .IN4(na350_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x94y69     80'h00_0018_00_0000_0888_77B3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1767_1 ( .OUT(na1767_1), .IN1(1'b0), .IN2(~na608_1), .IN3(na600_2), .IN4(~na102_2), .IN5(~na819_1), .IN6(~na2033_2), .IN7(~na1561_1),
                      .IN8(~na102_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x90y60     80'h00_0078_00_0000_0C88_C3CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1769_1 ( .OUT(na1769_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1770_1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1769_4 ( .OUT(na1769_2), .IN1(na913_2), .IN2(1'b1), .IN3(1'b1), .IN4(na49_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x77y74     80'h00_0018_00_0000_0888_77B3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1770_1 ( .OUT(na1770_1), .IN1(1'b0), .IN2(~na628_1), .IN3(na574_1), .IN4(~na102_2), .IN5(~na822_1), .IN6(~na2033_2), .IN7(~na1584_1),
                      .IN8(~na102_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x89y63     80'h00_0078_00_0000_0C88_C3CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1772_1 ( .OUT(na1772_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1773_1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1772_4 ( .OUT(na1772_2), .IN1(1'b1), .IN2(na567_1), .IN3(1'b1), .IN4(na1070_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x83y66     80'h00_0018_00_0000_0888_77B5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1773_1 ( .OUT(na1773_1), .IN1(~na635_1), .IN2(1'b0), .IN3(na556_1), .IN4(~na102_2), .IN5(~na1592_1), .IN6(~na1909_2), .IN7(~na825_1),
                      .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x85y64     80'h00_0018_00_0000_0888_7573
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1775_1 ( .OUT(na1775_1), .IN1(1'b0), .IN2(~na642_1), .IN3(~na1603_1), .IN4(~na102_1), .IN5(~na643_1), .IN6(1'b0), .IN7(~na828_1),
                      .IN8(~na1065_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y54     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1778_4 ( .OUT(na1778_2), .IN1(na1942_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1779_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y62     80'h00_0018_00_0000_0888_7755
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1779_1 ( .OUT(na1779_1), .IN1(~na648_1), .IN2(1'b0), .IN3(~na649_1), .IN4(1'b0), .IN5(~na831_1), .IN6(~na2033_2), .IN7(~na1612_1),
                      .IN8(~na102_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x92y61     80'h00_0078_00_0000_0C88_C3AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1782_1 ( .OUT(na1782_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1783_1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1782_4 ( .OUT(na1782_2), .IN1(na943_1), .IN2(1'b1), .IN3(na346_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x77y54     80'h00_0018_00_0000_0888_7753
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1783_1 ( .OUT(na1783_1), .IN1(1'b0), .IN2(~na664_1), .IN3(~na665_1), .IN4(1'b0), .IN5(~na836_1), .IN6(~na2033_2), .IN7(~na1631_1),
                      .IN8(~na102_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y64     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1788_4 ( .OUT(na1788_2), .IN1(1'b1), .IN2(na89_1), .IN3(1'b1), .IN4(~na418_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y55     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1790_4 ( .OUT(na1790_2), .IN1(na1942_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1791_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x80y60     80'h00_0018_00_0000_0888_FB73
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1791_1 ( .OUT(na1791_1), .IN1(1'b0), .IN2(~na845_1), .IN3(~na1389_1), .IN4(~na102_1), .IN5(na431_1), .IN6(~na101_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y60     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1793_1 ( .OUT(na1793_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na89_1), .IN7(na460_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y53     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1795_1 ( .OUT(na1795_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1796_1), .IN6(1'b1), .IN7(1'b1), .IN8(na350_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x83y65     80'h00_0018_00_0000_0888_FB75
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1796_1 ( .OUT(na1796_1), .IN1(~na848_1), .IN2(1'b0), .IN3(~na1420_1), .IN4(~na102_1), .IN5(na469_1), .IN6(~na101_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x59y128     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1797_4 ( .OUT(na1797_2), .IN1(1'b1), .IN2(1'b1), .IN3(na75_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1797_6 ( .RAM_O2(na1797_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1797_2), .COMP_OUT(1'b0) );
// C_///AND/      x61y128     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1798_4 ( .OUT(na1798_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na77_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1798_6 ( .RAM_O2(na1798_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1798_2), .COMP_OUT(1'b0) );
// C_///AND/      x65y128     80'h08_0060_00_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1799_4 ( .OUT(na1799_2), .IN1(1'b1), .IN2(~na146_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1799_6 ( .RAM_O2(na1799_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1799_2), .COMP_OUT(1'b0) );
// C_///AND/      x67y128     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1800_4 ( .OUT(na1800_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na151_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1800_6 ( .RAM_O2(na1800_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1800_2), .COMP_OUT(1'b0) );
// C_///AND/      x69y128     80'h08_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1801_4 ( .OUT(na1801_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na156_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1801_6 ( .RAM_O2(na1801_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1801_2), .COMP_OUT(1'b0) );
// C_///AND/      x73y128     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1802_4 ( .OUT(na1802_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na161_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1802_6 ( .RAM_O2(na1802_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1802_2), .COMP_OUT(1'b0) );
// C_///AND/      x75y128     80'h08_0060_00_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1803_4 ( .OUT(na1803_2), .IN1(1'b1), .IN2(~na166_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1803_6 ( .RAM_O2(na1803_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1803_2), .COMP_OUT(1'b0) );
// C_///AND/      x77y128     80'h08_0060_00_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1804_4 ( .OUT(na1804_2), .IN1(1'b1), .IN2(~na171_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1804_6 ( .RAM_O2(na1804_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1804_2), .COMP_OUT(1'b0) );
// C_///AND/      x81y128     80'h08_0060_00_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1805_4 ( .OUT(na1805_2), .IN1(~na176_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1805_6 ( .RAM_O2(na1805_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1805_2), .COMP_OUT(1'b0) );
// C_///AND/      x83y128     80'h08_0060_00_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1806_4 ( .OUT(na1806_2), .IN1(1'b1), .IN2(~na181_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1806_6 ( .RAM_O2(na1806_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1806_2), .COMP_OUT(1'b0) );
// C_///AND/      x87y128     80'h08_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1807_4 ( .OUT(na1807_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na186_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1807_6 ( .RAM_O2(na1807_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1807_2), .COMP_OUT(1'b0) );
// C_///AND/      x89y128     80'h08_0060_00_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1808_4 ( .OUT(na1808_2), .IN1(~na191_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1808_6 ( .RAM_O2(na1808_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1808_2), .COMP_OUT(1'b0) );
// C_///AND/      x91y128     80'h08_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1809_4 ( .OUT(na1809_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na106_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1809_6 ( .RAM_O2(na1809_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1809_2), .COMP_OUT(1'b0) );
// C_///AND/      x103y128     80'h08_0060_00_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1810_4 ( .OUT(na1810_2), .IN1(~na196_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1810_6 ( .RAM_O2(na1810_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1810_2), .COMP_OUT(1'b0) );
// C_///AND/      x105y128     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1811_4 ( .OUT(na1811_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na201_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1811_6 ( .RAM_O2(na1811_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1811_2), .COMP_OUT(1'b0) );
// C_///AND/      x107y128     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1812_4 ( .OUT(na1812_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na206_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1812_6 ( .RAM_O2(na1812_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1812_2), .COMP_OUT(1'b0) );
// C_///AND/      x111y128     80'h08_0060_00_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1813_4 ( .OUT(na1813_2), .IN1(~na211_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1813_6 ( .RAM_O2(na1813_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1813_2), .COMP_OUT(1'b0) );
// C_///AND/      x113y128     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1814_4 ( .OUT(na1814_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1814_6 ( .RAM_O2(na1814_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1814_2), .COMP_OUT(1'b0) );
// C_///AND/      x117y128     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1815_4 ( .OUT(na1815_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1815_6 ( .RAM_O2(na1815_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1815_2), .COMP_OUT(1'b0) );
// C_///AND/      x119y128     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1816_4 ( .OUT(na1816_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1816_6 ( .RAM_O2(na1816_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1816_2), .COMP_OUT(1'b0) );
// C_///AND/      x121y128     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1817_4 ( .OUT(na1817_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1817_6 ( .RAM_O2(na1817_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1817_2), .COMP_OUT(1'b0) );
// C_///AND/      x125y128     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1818_4 ( .OUT(na1818_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1818_6 ( .RAM_O2(na1818_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1818_2), .COMP_OUT(1'b0) );
// C_///AND/      x127y128     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1819_4 ( .OUT(na1819_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1819_6 ( .RAM_O2(na1819_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1819_2), .COMP_OUT(1'b0) );
// C_///AND/      x129y128     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1820_4 ( .OUT(na1820_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na111_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1820_6 ( .RAM_O2(na1820_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1820_2), .COMP_OUT(1'b0) );
// C_///AND/      x133y128     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1821_4 ( .OUT(na1821_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1821_6 ( .RAM_O2(na1821_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1821_2), .COMP_OUT(1'b0) );
// C_///AND/      x135y128     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1822_4 ( .OUT(na1822_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1822_6 ( .RAM_O2(na1822_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1822_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y27     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1823_4 ( .OUT(na1823_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na116_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1823_6 ( .RAM_O2(na1823_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1823_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y29     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1824_4 ( .OUT(na1824_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na121_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1824_6 ( .RAM_O2(na1824_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1824_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y31     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1825_4 ( .OUT(na1825_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na126_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1825_6 ( .RAM_O2(na1825_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1825_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y35     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1826_4 ( .OUT(na1826_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na131_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1826_6 ( .RAM_O2(na1826_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1826_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y37     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1827_4 ( .OUT(na1827_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na136_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1827_6 ( .RAM_O2(na1827_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1827_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y39     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1828_4 ( .OUT(na1828_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na141_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1828_6 ( .RAM_O2(na1828_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1828_2), .COMP_OUT(1'b0) );
// C_///AND/      x101y1     80'h08_0060_00_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1829_4 ( .OUT(na1829_2), .IN1(1'b1), .IN2(~na736_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1829_6 ( .RAM_O2(na1829_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1829_2), .COMP_OUT(1'b0) );
// C_///AND/      x107y1     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1830_4 ( .OUT(na1830_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1302_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1830_6 ( .RAM_O2(na1830_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1830_2), .COMP_OUT(1'b0) );
// C_///AND/      x109y1     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1831_4 ( .OUT(na1831_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1301_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1831_6 ( .RAM_O2(na1831_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1831_2), .COMP_OUT(1'b0) );
// C_///AND/      x113y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1832_4 ( .OUT(na1832_2), .IN1(1'b1), .IN2(na218_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1832_6 ( .RAM_O2(na1832_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1832_2), .COMP_OUT(1'b0) );
// C_///AND/      x115y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1833_4 ( .OUT(na1833_2), .IN1(1'b1), .IN2(na219_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1833_6 ( .RAM_O2(na1833_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1833_2), .COMP_OUT(1'b0) );
// C_///AND/      x117y1     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1834_4 ( .OUT(na1834_2), .IN1(na220_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1834_6 ( .RAM_O2(na1834_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1834_2), .COMP_OUT(1'b0) );
// C_///AND/      x121y1     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1835_4 ( .OUT(na1835_2), .IN1(na221_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1835_6 ( .RAM_O2(na1835_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1835_2), .COMP_OUT(1'b0) );
// C_///AND/      x123y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1836_4 ( .OUT(na1836_2), .IN1(1'b1), .IN2(na222_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1836_6 ( .RAM_O2(na1836_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1836_2), .COMP_OUT(1'b0) );
// C_///AND/      x125y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1837_4 ( .OUT(na1837_2), .IN1(1'b1), .IN2(na223_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1837_6 ( .RAM_O2(na1837_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1837_2), .COMP_OUT(1'b0) );
// C_///AND/      x129y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1838_4 ( .OUT(na1838_2), .IN1(1'b1), .IN2(na224_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1838_6 ( .RAM_O2(na1838_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1838_2), .COMP_OUT(1'b0) );
// C_///AND/      x131y1     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1839_4 ( .OUT(na1839_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na225_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1839_6 ( .RAM_O2(na1839_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1839_2), .COMP_OUT(1'b0) );
// C_///AND/      x133y1     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1840_4 ( .OUT(na1840_2), .IN1(1'b1), .IN2(1'b1), .IN3(na226_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1840_6 ( .RAM_O2(na1840_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1840_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y25     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1841_4 ( .OUT(na1841_2), .IN1(1'b1), .IN2(1'b1), .IN3(na227_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1841_6 ( .RAM_O2(na1841_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1841_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y27     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1842_4 ( .OUT(na1842_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1299_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1842_6 ( .RAM_O2(na1842_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1842_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y31     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1843_4 ( .OUT(na1843_2), .IN1(1'b1), .IN2(1'b1), .IN3(na228_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1843_6 ( .RAM_O2(na1843_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1843_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y33     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1844_4 ( .OUT(na1844_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na229_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1844_6 ( .RAM_O2(na1844_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1844_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y35     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1845_4 ( .OUT(na1845_2), .IN1(1'b1), .IN2(1'b1), .IN3(na230_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1845_6 ( .RAM_O2(na1845_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1845_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y39     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1846_4 ( .OUT(na1846_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na231_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1846_6 ( .RAM_O2(na1846_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1846_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y41     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1847_4 ( .OUT(na1847_2), .IN1(na232_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1847_6 ( .RAM_O2(na1847_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1847_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y43     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1848_4 ( .OUT(na1848_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na233_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1848_6 ( .RAM_O2(na1848_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1848_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y47     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1849_4 ( .OUT(na1849_2), .IN1(1'b1), .IN2(na234_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1849_6 ( .RAM_O2(na1849_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1849_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y49     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1850_4 ( .OUT(na1850_2), .IN1(na235_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1850_6 ( .RAM_O2(na1850_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1850_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y53     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1851_4 ( .OUT(na1851_2), .IN1(1'b1), .IN2(1'b1), .IN3(na236_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1851_6 ( .RAM_O2(na1851_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1851_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y55     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1852_4 ( .OUT(na1852_2), .IN1(na237_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1852_6 ( .RAM_O2(na1852_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1852_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y57     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1853_4 ( .OUT(na1853_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1298_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1853_6 ( .RAM_O2(na1853_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1853_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y69     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1854_4 ( .OUT(na1854_2), .IN1(na238_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1854_6 ( .RAM_O2(na1854_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1854_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y71     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1855_4 ( .OUT(na1855_2), .IN1(1'b1), .IN2(na239_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1855_6 ( .RAM_O2(na1855_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1855_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y73     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1856_4 ( .OUT(na1856_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1297_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1856_6 ( .RAM_O2(na1856_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1856_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y77     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1857_4 ( .OUT(na1857_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1295_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1857_6 ( .RAM_O2(na1857_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1857_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y79     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1858_4 ( .OUT(na1858_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1294_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1858_6 ( .RAM_O2(na1858_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1858_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y83     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1859_4 ( .OUT(na1859_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1293_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1859_6 ( .RAM_O2(na1859_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1859_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y85     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1860_4 ( .OUT(na1860_2), .IN1(na216_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1860_6 ( .RAM_O2(na1860_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1860_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y87     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1861_4 ( .OUT(na1861_2), .IN1(na217_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1861_6 ( .RAM_O2(na1861_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1861_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y91     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1862_4 ( .OUT(na1862_2), .IN1(na737_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1862_6 ( .RAM_O2(na1862_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1862_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y93     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1863_4 ( .OUT(na1863_2), .IN1(na739_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1863_6 ( .RAM_O2(na1863_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1863_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y95     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1864_4 ( .OUT(na1864_2), .IN1(1'b1), .IN2(na740_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1864_6 ( .RAM_O2(na1864_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1864_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y89     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1865_4 ( .OUT(na1865_2), .IN1(na741_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1865_6 ( .RAM_O2(na1865_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1865_2), .COMP_OUT(1'b0) );
// C_////Bridge      x92y69     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1866_5 ( .OUT(na1866_2), .IN1(na3_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1867_5 ( .OUT(na1867_2), .IN1(1'b0), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y66     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1868_5 ( .OUT(na1868_2), .IN1(1'b0), .IN2(na4_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1869_5 ( .OUT(na1869_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y60     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1870_5 ( .OUT(na1870_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na5_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y76     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1871_5 ( .OUT(na1871_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na7_1) );
// C_////Bridge      x90y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1872_5 ( .OUT(na1872_2), .IN1(1'b0), .IN2(na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y78     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1873_5 ( .OUT(na1873_2), .IN1(1'b0), .IN2(na8_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y66     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1874_5 ( .OUT(na1874_2), .IN1(1'b0), .IN2(na9_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y75     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1875_5 ( .OUT(na1875_2), .IN1(1'b0), .IN2(1'b0), .IN3(na10_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y74     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1876_5 ( .OUT(na1876_2), .IN1(1'b0), .IN2(1'b0), .IN3(na10_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y66     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1877_5 ( .OUT(na1877_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na11_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y58     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1878_5 ( .OUT(na1878_2), .IN1(1'b0), .IN2(na12_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y50     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1879_5 ( .OUT(na1879_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na13_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y47     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1880_5 ( .OUT(na1880_2), .IN1(na14_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y61     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1881_5 ( .OUT(na1881_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na15_1) );
// C_////Bridge      x80y52     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1882_5 ( .OUT(na1882_2), .IN1(1'b0), .IN2(na16_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y52     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1883_5 ( .OUT(na1883_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na17_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y54     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1884_5 ( .OUT(na1884_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na18_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y48     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1885_5 ( .OUT(na1885_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na19_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y64     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1886_5 ( .OUT(na1886_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na20_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y54     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1887_5 ( .OUT(na1887_2), .IN1(na23_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y68     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1888_5 ( .OUT(na1888_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na24_1) );
// C_////Bridge      x74y54     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1889_5 ( .OUT(na1889_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na25_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y56     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1890_5 ( .OUT(na1890_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na26_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y70     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1891_5 ( .OUT(na1891_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na28_1) );
// C_////Bridge      x84y52     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1892_5 ( .OUT(na1892_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na30_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y72     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1893_5 ( .OUT(na1893_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na31_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y50     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1894_5 ( .OUT(na1894_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na33_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y48     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1895_5 ( .OUT(na1895_2), .IN1(na35_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y74     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1896_5 ( .OUT(na1896_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na36_1) );
// C_////Bridge      x74y52     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1897_5 ( .OUT(na1897_2), .IN1(1'b0), .IN2(na37_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y59     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1898_5 ( .OUT(na1898_2), .IN1(na38_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y70     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1899_5 ( .OUT(na1899_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na44_2) );
// C_////Bridge      x91y62     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1900_5 ( .OUT(na1900_2), .IN1(na45_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y67     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1901_5 ( .OUT(na1901_2), .IN1(na45_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y68     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1902_5 ( .OUT(na1902_2), .IN1(na45_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y63     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1903_5 ( .OUT(na1903_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na49_1) );
// C_////Bridge      x81y52     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1904_5 ( .OUT(na1904_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na83_2), .IN8(1'b0) );
// C_////Bridge      x84y69     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1905_5 ( .OUT(na1905_2), .IN1(na84_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y60     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1906_5 ( .OUT(na1906_2), .IN1(na84_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y66     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1907_5 ( .OUT(na1907_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na101_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y65     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1908_5 ( .OUT(na1908_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na102_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y64     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1909_5 ( .OUT(na1909_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na102_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y61     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1910_5 ( .OUT(na1910_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na102_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y68     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1911_5 ( .OUT(na1911_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na102_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y61     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1912_5 ( .OUT(na1912_2), .IN1(1'b0), .IN2(1'b0), .IN3(na247_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1913_5 ( .OUT(na1913_2), .IN1(1'b0), .IN2(1'b0), .IN3(na247_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y55     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1914_5 ( .OUT(na1914_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na249_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y56     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1915_5 ( .OUT(na1915_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na250_1) );
// C_////Bridge      x95y72     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1916_5 ( .OUT(na1916_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na250_2) );
// C_////Bridge      x92y64     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1917_5 ( .OUT(na1917_2), .IN1(1'b0), .IN2(na258_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y62     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1918_5 ( .OUT(na1918_2), .IN1(1'b0), .IN2(na258_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y58     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1919_5 ( .OUT(na1919_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na260_1) );
// C_////Bridge      x85y80     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1920_5 ( .OUT(na1920_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na260_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y68     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1921_5 ( .OUT(na1921_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na262_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y66     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1922_5 ( .OUT(na1922_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na262_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y70     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1923_5 ( .OUT(na1923_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na264_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y68     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1924_5 ( .OUT(na1924_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na264_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y70     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1925_5 ( .OUT(na1925_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na266_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y74     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1926_5 ( .OUT(na1926_2), .IN1(1'b0), .IN2(na266_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y76     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1927_5 ( .OUT(na1927_2), .IN1(1'b0), .IN2(na268_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y72     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1928_5 ( .OUT(na1928_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na268_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y76     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1929_5 ( .OUT(na1929_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na269_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y76     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1930_5 ( .OUT(na1930_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na273_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y72     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1931_5 ( .OUT(na1931_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na284_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y64     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1932_5 ( .OUT(na1932_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na298_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y70     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1933_5 ( .OUT(na1933_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na303_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1934_5 ( .OUT(na1934_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na307_1) );
// C_////Bridge      x77y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1935_5 ( .OUT(na1935_2), .IN1(na311_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y80     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1936_5 ( .OUT(na1936_2), .IN1(1'b0), .IN2(na322_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y69     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1937_5 ( .OUT(na1937_2), .IN1(1'b0), .IN2(1'b0), .IN3(na326_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1938_5 ( .OUT(na1938_2), .IN1(1'b0), .IN2(1'b0), .IN3(na327_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1939_5 ( .OUT(na1939_2), .IN1(1'b0), .IN2(1'b0), .IN3(na327_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y60     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1940_5 ( .OUT(na1940_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na335_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1941_5 ( .OUT(na1941_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na350_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1942_5 ( .OUT(na1942_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na350_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y56     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1943_5 ( .OUT(na1943_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na350_2) );
// C_////Bridge      x84y66     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1944_5 ( .OUT(na1944_2), .IN1(1'b0), .IN2(na356_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1945_5 ( .OUT(na1945_2), .IN1(na359_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1946_5 ( .OUT(na1946_2), .IN1(1'b0), .IN2(1'b0), .IN3(na361_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y81     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1947_5 ( .OUT(na1947_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na363_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y78     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1948_5 ( .OUT(na1948_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na370_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y69     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1949_5 ( .OUT(na1949_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na378_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y80     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1950_5 ( .OUT(na1950_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na396_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1951_5 ( .OUT(na1951_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na402_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y66     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1952_5 ( .OUT(na1952_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na410_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y78     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1953_5 ( .OUT(na1953_2), .IN1(1'b0), .IN2(na430_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y78     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1954_5 ( .OUT(na1954_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na465_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y76     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1955_5 ( .OUT(na1955_2), .IN1(1'b0), .IN2(na468_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1956_5 ( .OUT(na1956_2), .IN1(1'b0), .IN2(1'b0), .IN3(na470_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y61     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1957_5 ( .OUT(na1957_2), .IN1(1'b0), .IN2(1'b0), .IN3(na479_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y53     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1958_5 ( .OUT(na1958_2), .IN1(na496_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y48     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1959_5 ( .OUT(na1959_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na509_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y49     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1960_5 ( .OUT(na1960_2), .IN1(1'b0), .IN2(1'b0), .IN3(na510_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y59     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1961_5 ( .OUT(na1961_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na525_1), .IN8(1'b0) );
// C_////Bridge      x91y76     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1962_5 ( .OUT(na1962_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na538_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y63     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1963_5 ( .OUT(na1963_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na556_1), .IN8(1'b0) );
// C_////Bridge      x83y57     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1964_5 ( .OUT(na1964_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na567_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y69     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1965_5 ( .OUT(na1965_2), .IN1(1'b0), .IN2(1'b0), .IN3(na574_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y51     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1966_5 ( .OUT(na1966_2), .IN1(1'b0), .IN2(1'b0), .IN3(na600_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y75     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1967_5 ( .OUT(na1967_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na777_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y53     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1968_5 ( .OUT(na1968_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na870_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y53     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1969_5 ( .OUT(na1969_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na875_1) );
// C_////Bridge      x75y50     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1970_5 ( .OUT(na1970_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na883_1), .IN8(1'b0) );
// C_////Bridge      x81y77     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1971_5 ( .OUT(na1971_2), .IN1(1'b0), .IN2(1'b0), .IN3(na885_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y79     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1972_5 ( .OUT(na1972_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na885_2), .IN8(1'b0) );
// C_////Bridge      x83y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1973_5 ( .OUT(na1973_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na887_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1974_5 ( .OUT(na1974_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na887_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y83     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1975_5 ( .OUT(na1975_2), .IN1(1'b0), .IN2(1'b0), .IN3(na889_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y75     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1976_5 ( .OUT(na1976_2), .IN1(1'b0), .IN2(1'b0), .IN3(na889_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y81     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1977_5 ( .OUT(na1977_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na891_1) );
// C_////Bridge      x93y79     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1978_5 ( .OUT(na1978_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na891_2) );
// C_////Bridge      x79y83     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1979_5 ( .OUT(na1979_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na893_1), .IN8(1'b0) );
// C_////Bridge      x87y83     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1980_5 ( .OUT(na1980_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na893_2), .IN8(1'b0) );
// C_////Bridge      x77y57     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1981_5 ( .OUT(na1981_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na894_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y56     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1982_5 ( .OUT(na1982_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na894_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1983_5 ( .OUT(na1983_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na896_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1984_5 ( .OUT(na1984_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na896_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y77     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1985_5 ( .OUT(na1985_2), .IN1(1'b0), .IN2(1'b0), .IN3(na898_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y75     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1986_5 ( .OUT(na1986_2), .IN1(1'b0), .IN2(1'b0), .IN3(na899_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y71     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1987_5 ( .OUT(na1987_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na900_1) );
// C_////Bridge      x97y71     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1988_5 ( .OUT(na1988_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na901_1), .IN8(1'b0) );
// C_////Bridge      x99y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1989_5 ( .OUT(na1989_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na902_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y71     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1990_5 ( .OUT(na1990_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na902_2) );
// C_////Bridge      x99y71     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1991_5 ( .OUT(na1991_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na904_1), .IN8(1'b0) );
// C_////Bridge      x101y73     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1992_5 ( .OUT(na1992_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na904_2), .IN8(1'b0) );
// C_////Bridge      x97y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1993_5 ( .OUT(na1993_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na906_1) );
// C_////Bridge      x91y73     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1994_5 ( .OUT(na1994_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na906_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y72     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1995_5 ( .OUT(na1995_2), .IN1(na909_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y72     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1996_5 ( .OUT(na1996_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na913_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y76     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1997_5 ( .OUT(na1997_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na917_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1998_5 ( .OUT(na1998_2), .IN1(1'b0), .IN2(na931_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y67     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1999_5 ( .OUT(na1999_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na935_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y73     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2000_5 ( .OUT(na2000_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na939_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y61     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2001_5 ( .OUT(na2001_2), .IN1(1'b0), .IN2(na944_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y61     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2002_5 ( .OUT(na2002_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na984_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y56     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2003_5 ( .OUT(na2003_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na985_1), .IN8(1'b0) );
// C_////Bridge      x65y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2004_5 ( .OUT(na2004_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na987_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y68     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2005_5 ( .OUT(na2005_2), .IN1(1'b0), .IN2(1'b0), .IN3(na989_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y57     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2006_5 ( .OUT(na2006_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na991_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y60     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2007_5 ( .OUT(na2007_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na993_1), .IN8(1'b0) );
// C_////Bridge      x65y61     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2008_5 ( .OUT(na2008_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na996_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y60     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2009_5 ( .OUT(na2009_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na998_1), .IN8(1'b0) );
// C_////Bridge      x65y65     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2010_5 ( .OUT(na2010_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1000_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y68     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2011_5 ( .OUT(na2011_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1002_1), .IN8(1'b0) );
// C_////Bridge      x71y57     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2012_5 ( .OUT(na2012_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1004_1) );
// C_////Bridge      x73y56     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2013_5 ( .OUT(na2013_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1006_1), .IN8(1'b0) );
// C_////Bridge      x71y58     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2014_5 ( .OUT(na2014_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1007_1), .IN8(1'b0) );
// C_////Bridge      x75y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2015_5 ( .OUT(na2015_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1011_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y62     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2016_5 ( .OUT(na2016_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1013_1), .IN8(1'b0) );
// C_////Bridge      x71y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2017_5 ( .OUT(na2017_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1015_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y61     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2018_5 ( .OUT(na2018_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1023_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y59     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2019_5 ( .OUT(na2019_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1055_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2020_5 ( .OUT(na2020_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1055_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y54     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2021_5 ( .OUT(na2021_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1056_1) );
// C_////Bridge      x79y52     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2022_5 ( .OUT(na2022_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1058_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y59     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2023_5 ( .OUT(na2023_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1058_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y67     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2024_5 ( .OUT(na2024_2), .IN1(na1059_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2025_5 ( .OUT(na2025_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1060_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y50     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2026_5 ( .OUT(na2026_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1061_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y69     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2027_5 ( .OUT(na2027_2), .IN1(na1061_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y59     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2028_5 ( .OUT(na2028_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1062_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y51     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2029_5 ( .OUT(na2029_2), .IN1(1'b0), .IN2(na1063_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y62     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2030_5 ( .OUT(na2030_2), .IN1(1'b0), .IN2(na1063_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y49     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2031_5 ( .OUT(na2031_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1064_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y53     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2032_5 ( .OUT(na2032_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1065_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y58     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2033_5 ( .OUT(na2033_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1065_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y66     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2034_5 ( .OUT(na2034_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1066_1) );
// C_////Bridge      x91y68     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2035_5 ( .OUT(na2035_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1067_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y68     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2036_5 ( .OUT(na2036_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1068_2) );
// C_////Bridge      x91y72     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2037_5 ( .OUT(na2037_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1069_2) );
// C_////Bridge      x93y70     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2038_5 ( .OUT(na2038_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1070_1) );
// C_////Bridge      x82y63     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2039_5 ( .OUT(na2039_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1077_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y57     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2040_5 ( .OUT(na2040_2), .IN1(na1077_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y56     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2041_5 ( .OUT(na2041_2), .IN1(na1077_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y63     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2042_5 ( .OUT(na2042_2), .IN1(na1079_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y57     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2043_5 ( .OUT(na2043_2), .IN1(na1079_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x84y59     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2044_5 ( .OUT(na2044_2), .IN1(na1081_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y59     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2045_5 ( .OUT(na2045_2), .IN1(na1081_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y74     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2046_5 ( .OUT(na2046_2), .IN1(1'b0), .IN2(na1228_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2047_5 ( .OUT(na2047_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1277_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y50     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2048_5 ( .OUT(na2048_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1277_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y45     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2049_5 ( .OUT(na2049_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1278_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y51     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2050_5 ( .OUT(na2050_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1279_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y52     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2051_5 ( .OUT(na2051_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1281_1), .IN8(1'b0) );
// C_////Bridge      x81y48     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2052_5 ( .OUT(na2052_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1282_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y45     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2053_5 ( .OUT(na2053_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1283_1) );
// C_////Bridge      x81y45     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2054_5 ( .OUT(na2054_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1285_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y66     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2055_5 ( .OUT(na2055_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1285_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y71     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2056_5 ( .OUT(na2056_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1286_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y48     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2057_5 ( .OUT(na2057_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1286_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y44     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2058_5 ( .OUT(na2058_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1287_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y45     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2059_5 ( .OUT(na2059_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1289_1) );
// C_////Bridge      x61y61     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2060_5 ( .OUT(na2060_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1290_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2061_5 ( .OUT(na2061_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1291_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2062_5 ( .OUT(na2062_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1306_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x76y74     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2063_5 ( .OUT(na2063_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1307_1), .IN8(1'b0) );
// C_////Bridge      x61y65     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2064_5 ( .OUT(na2064_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1310_1) );
// C_////Bridge      x62y66     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2065_5 ( .OUT(na2065_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1311_2), .IN8(1'b0) );
// C_////Bridge      x73y67     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2066_5 ( .OUT(na2066_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1313_1), .IN8(1'b0) );
// C_////Bridge      x67y52     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2067_5 ( .OUT(na2067_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1314_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x69y54     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2068_5 ( .OUT(na2068_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1315_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y51     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2069_5 ( .OUT(na2069_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1317_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2070_5 ( .OUT(na2070_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1317_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y47     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2071_5 ( .OUT(na2071_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1318_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y66     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2072_5 ( .OUT(na2072_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1318_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y77     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2073_5 ( .OUT(na2073_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1332_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2074_5 ( .OUT(na2074_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1337_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y62     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2075_5 ( .OUT(na2075_2), .IN1(na1341_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y50     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2076_5 ( .OUT(na2076_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1341_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y75     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2077_5 ( .OUT(na2077_2), .IN1(1'b0), .IN2(na1350_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y47     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2078_5 ( .OUT(na2078_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1359_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y65     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2079_5 ( .OUT(na2079_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1372_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y43     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2080_5 ( .OUT(na2080_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1393_1) );
// C_////Bridge      x85y61     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2081_5 ( .OUT(na2081_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1399_1), .IN8(1'b0) );
// C_////Bridge      x95y47     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2082_5 ( .OUT(na2082_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1410_1) );
// C_////Bridge      x79y75     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2083_5 ( .OUT(na2083_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1418_1), .IN8(1'b0) );
// C_////Bridge      x97y45     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2084_5 ( .OUT(na2084_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1424_1) );
// C_////Bridge      x73y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2085_5 ( .OUT(na2085_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1430_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y53     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2086_5 ( .OUT(na2086_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1433_1) );
// C_////Bridge      x73y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2087_5 ( .OUT(na2087_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1436_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y45     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2088_5 ( .OUT(na2088_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1437_1) );
// C_////Bridge      x71y51     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2089_5 ( .OUT(na2089_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1442_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y49     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2090_5 ( .OUT(na2090_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1454_2), .IN8(1'b0) );
// C_////Bridge      x71y49     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2091_5 ( .OUT(na2091_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1455_1), .IN8(1'b0) );
// C_////Bridge      x77y55     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2092_5 ( .OUT(na2092_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1459_2) );
// C_////Bridge      x81y51     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2093_5 ( .OUT(na2093_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1463_1) );
// C_////Bridge      x77y49     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2094_5 ( .OUT(na2094_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1468_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y49     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2095_5 ( .OUT(na2095_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1474_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y48     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2096_5 ( .OUT(na2096_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1475_2) );
// C_////Bridge      x79y50     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2097_5 ( .OUT(na2097_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1478_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y58     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2098_5 ( .OUT(na2098_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1480_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y67     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2099_5 ( .OUT(na2099_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1481_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x75y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2100_5 ( .OUT(na2100_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1484_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y58     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2101_5 ( .OUT(na2101_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1491_2) );
// C_////Bridge      x75y58     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2102_5 ( .OUT(na2102_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1492_1) );
// C_////Bridge      x73y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2103_5 ( .OUT(na2103_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1493_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2104_5 ( .OUT(na2104_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1493_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y65     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2105_5 ( .OUT(na2105_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1494_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y60     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2106_5 ( .OUT(na2106_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1496_1), .IN8(1'b0) );
// C_////Bridge      x63y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2107_5 ( .OUT(na2107_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1497_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y51     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2108_5 ( .OUT(na2108_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1503_1) );
// C_////Bridge      x87y63     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2109_5 ( .OUT(na2109_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1504_2), .IN8(1'b0) );
// C_////Bridge      x73y47     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2110_5 ( .OUT(na2110_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1509_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y49     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2111_5 ( .OUT(na2111_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1514_1) );
// C_////Bridge      x79y47     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2112_5 ( .OUT(na2112_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1517_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y51     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2113_5 ( .OUT(na2113_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1518_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y47     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2114_5 ( .OUT(na2114_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1520_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y58     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2115_5 ( .OUT(na2115_2), .IN1(1'b0), .IN2(na1568_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y60     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a2116_5 ( .OUT(na2116_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1782_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
endmodule
