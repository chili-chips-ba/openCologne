serdes_inst: CC_SERDES
generic map (
  CCAG_CFG_PARAM           => "", // legacy
  SERDES_ENABLE            => 0,

  TX_SEL_PRE               => 0,
  TX_SEL_POST              => 0,
  TX_AMP                   => 15,
  TX_BRANCH_EN_PRE         => 0,
  TX_BRANCH_EN_MAIN        => X"3F",
  TX_BRANCH_EN_POST        => 0,
  TX_TAIL_CASCODE          => 4,
  TX_DC_ENABLE             => 63,
  TX_DC_OFFSET             => 0,
  TX_CM_RAISE              => 0,
  TX_CM_THRESHOLD_0        => 14,
  TX_CM_THRESHOLD_1        => 16,
  TX_SEL_PRE_EI            => 0,
  TX_SEL_POST_EI           => 0,
  TX_AMP_EI                => 15,
  TX_BRANCH_EN_PRE_EI      => 0,
  TX_BRANCH_EN_MAIN_EI     => X"3F",
  TX_BRANCH_EN_POST_EI     => 0,
  TX_TAIL_CASCODE_EI       => 4,
  TX_DC_ENABLE_EI          => 63,
  TX_DC_OFFSET_EI          => 0,
  TX_CM_RAISE_EI           => 0,
  TX_CM_THRESHOLD_0_EI     => 14,
  TX_CM_THRESHOLD_1_EI     => 16,
  TX_SEL_PRE_RXDET         => 0,
  TX_SEL_POST_RXDET        => 0,
  TX_AMP_RXDET             => 15,
  TX_BRANCH_EN_PRE_RXDET   => 0,
  TX_BRANCH_EN_MAIN_RXDET  => X"3F",
  TX_BRANCH_EN_POST_RXDET  => 0,
  TX_TAIL_CASCODE_RXDET    => 4,
  TX_DC_ENABLE_RXDET       => 63,
  TX_DC_OFFSET_RXDET       => 0,
  TX_CM_RAISE_RXDET        => 0,
  TX_CM_THRESHOLD_0_RXDET  => 14,
  TX_CM_THRESHOLD_1_RXDET  => 16,
  TX_CALIB_EN              => 0,
  TX_CALIB_OVR             => 0,
  TX_CALIB_VAL             => 0,
  TX_CM_REG_KI             => X"80",
  TX_CM_SAR_EN             => 0,
  TX_CM_REG_EN             => 1,
  TX_PMA_RESET_TIME        => 3,
  TX_PCS_RESET_TIME        => 3,
  TX_PCS_RESET_OVR         => 0,
  TX_PCS_RESET             => 0,
  TX_PMA_RESET_OVR         => 0,
  TX_PMA_RESET             => 0,
  TX_RESET_OVR             => 0,
  TX_RESET                 => 0,
  TX_PMA_LOOPBACK          => 0,
  TX_PCS_LOOPBACK          => 0,
  TX_DATAPATH_SEL          => 3,
  TX_PRBS_OVR              => 0,
  TX_PRBS_SEL              => 0,
  TX_PRBS_FORCE_ERR        => 0,
  TX_LOOPBACK_OVR          => 0,
  TX_POWERDOWN_OVR         => 0,
  TX_POWERDOWN_N           => 0,
  TX_ELEC_IDLE_OVR         => 0,
  TX_ELEC_IDLE             => 0,
  TX_DETECT_RX_OVR         => 0,
  TX_DETECT_RX             => 0,
  TX_POLARITY_OVR          => 0,
  TX_POLARITY              => 0,
  TX_8B10B_EN_OVR          => 0,
  TX_8B10B_EN              => 0,
  TX_DATA_OVR              => 0,
  TX_DATA_CNT              => 0,
  TX_DATA_VALID            => 0,

  RX_BUF_RESET_TIME        => 3,
  RX_PCS_RESET_TIME        => 3,
  RX_RESET_TIMER_PRESC     => 0,
  RX_RESETDONE_GATE        => 0,
  RX_CDR_RESET_TIME        => 3,
  RX_EQA_RESET_TIME        => 3,
  RX_PMA_RESET_TIME        => 3,
  RX_WAIT_CDR_LOCK         => 1,
  RX_CALIB_EN              => 0,
  RX_CALIB_OVR             => 0,
  RX_CALIB_VAL             => 0,
  RX_RTERM_VCMSEL          => 4,
  RX_RTERM_PD              => 0,
  RX_EQA_CKP_LF            => X"A3",
  RX_EQA_CKP_HF            => X"A3",
  RX_EQA_CKP_OFFSET        => X"01",
  RX_EN_EQA                => 0,
  RX_EQA_LOCK_CFG          => 0,
  RX_TH_MON1               => 8,
  RX_EN_EQA_EXT_VALUE      => 0,
  RX_TH_MON2               => 8,
  RX_TAPW                  => 8,
  RX_AFE_OFFSET            => 8,
  RX_EQA_CONFIG            => X"01C0",
  RX_AFE_PEAK              => 16,
  RX_AFE_GAIN              => 8,
  RX_AFE_VCMSEL            => 4,
  RX_CDR_CKP               => X"F8",
  RX_CDR_CKI               => 0,
  RX_CDR_TRANS_TH          => 128,
  RX_CDR_LOCK_CFG          => X"0B",
  RX_CDR_FREQ_ACC          => 0,
  RX_CDR_PHASE_ACC         => 0,
  RX_CDR_SET_ACC_CONFIG    => 0,
  RX_CDR_FORCE_LOCK        => 0,
  RX_ALIGN_MCOMMA_VALUE    => X"283",
  RX_MCOMMA_ALIGN_OVR      => 0,
  RX_MCOMMA_ALIGN          => 0,
  RX_ALIGN_PCOMMA_VALUE    => X"17C",
  RX_PCOMMA_ALIGN_OVR      => 0,
  RX_PCOMMA_ALIGN          => 0,
  RX_ALIGN_COMMA_WORD      => 0,
  RX_ALIGN_COMMA_ENABLE    => X"3FF",
  RX_SLIDE_MODE            => 0,
  RX_COMMA_DETECT_EN_OVR   => 0,
  RX_COMMA_DETECT_EN       => 0,
  RX_SLIDE                 => 0,
  RX_EYE_MEAS_EN           => 0,
  RX_EYE_MEAS_CFG          => 0,
  RX_MON_PH_OFFSET         => 0,
  RX_EI_BIAS               => 0,
  RX_EI_BW_SEL             => 4,
  RX_EN_EI_DETECTOR_OVR    => 0,
  RX_EN_EI_DETECTOR        => 0,
  RX_DATA_SEL              => 0,
  RX_BUF_BYPASS            => 0,
  RX_CLKCOR_USE            => 0,
  RX_CLKCOR_MIN_LAT        => 32,
  RX_CLKCOR_MAX_LAT        => 39,
  RX_CLKCOR_SEQ_1_0        => X"1F7",
  RX_CLKCOR_SEQ_1_1        => X"1F7",
  RX_CLKCOR_SEQ_1_2        => X"1F7",
  RX_CLKCOR_SEQ_1_3        => X"1F7",
  RX_PMA_LOOPBACK          => 0,
  RX_PCS_LOOPBACK          => 0,
  RX_DATAPATH_SEL          => 3,
  RX_PRBS_OVR              => 0,
  RX_PRBS_SEL              => 0,
  RX_LOOPBACK_OVR          => 0,
  RX_PRBS_CNT_RESET        => 0,
  RX_POWERDOWN_OVR         => 0,
  RX_POWERDOWN_N           => 0,
  RX_RESET_OVR             => 0,
  RX_RESET                 => 0,
  RX_PMA_RESET_OVR         => 0,
  RX_PMA_RESET             => 0,
  RX_EQA_RESET_OVR         => 0,
  RX_EQA_RESET             => 0,
  RX_CDR_RESET_OVR         => 0,
  RX_CDR_RESET             => 0,
  RX_PCS_RESET_OVR         => 0,
  RX_PCS_RESET             => 0,
  RX_BUF_RESET_OVR         => 0,
  RX_BUF_RESET             => 0,
  RX_POLARITY_OVR          => 0,
  RX_POLARITY              => 0,
  RX_8B10B_EN_OVR          => 0,
  RX_8B10B_EN              => 0,
  RX_8B10B_BYPASS          => 0,
  RX_BYTE_REALIGN          => 0,
  RX_DBG_EN                => 0,
  RX_DBG_SEL               => 0,
  RX_DBG_MODE              => 0,
  RX_DBG_SRAM_DELAY        => X"05",
  RX_DBG_ADDR              => 0,
  RX_DBG_RE                => 0,
  RX_DBG_WE                => 0,
  RX_DBG_DATA              => 0,

  PLL_EN_ADPLL_CTRL        => 0,
  PLL_CONFIG_SEL           => 0,
  PLL_SET_OP_LOCK          => 0,
  PLL_ENFORCE_LOCK         => 0,
  PLL_DISABLE_LOCK         => 0,
  PLL_LOCK_WINDOW          => 1,
  PLL_FAST_LOCK            => 1,
  PLL_SYNC_BYPASS          => 0,
  PLL_PFD_SELECT           => 0,
  PLL_REF_BYPASS           => 0,
  PLL_REF_SEL              => 0,
  PLL_REF_RTERM            => 1,
  PLL_FCNTRL               => 58,
  PLL_MAIN_DIVSEL          => 27,
  PLL_OUT_DIVSEL           => 0,
  PLL_CI                   => 3,
  PLL_CP                   => 80,
  PLL_AO                   => 0,
  PLL_SCAP                 => 0,
  PLL_FILTER_SHIFT         => 2,
  PLL_SAR_LIMIT            => 2,
  PLL_FT                   => 512,
  PLL_OPEN_LOOP            => 0,
  PLL_SCAP_AUTO_CAL        => 1,
  PLL_BISC_MODE            => 4,
  PLL_BISC_TIMER_MAX       => 15,
  PLL_BISC_OPT_DET_IND     => 0,
  PLL_BISC_PFD_SEL         => 0,
  PLL_BISC_DLY_DIR         => 0,
  PLL_BISC_COR_DLY         => 1,
  PLL_BISC_CAL_SIGN        => 0,
  PLL_BISC_CAL_AUTO        => 1,
  PLL_BISC_CP_MIN          => 4,
  PLL_BISC_CP_MAX          => 18,
  PLL_BISC_CP_START        => 12,
  PLL_BISC_DLY_PFD_MON_REF => 0,
  PLL_BISC_DLY_PFD_MON_DIV => 2
)
port map (
  TX_RESET_I             => TX_RESET_I,
  TX_PCS_RESET_I         => TX_PCS_RESET_I,
  TX_PMA_RESET_I         => TX_PMA_RESET_I,
  TX_POWER_DOWN_N_I      => TX_POWER_DOWN_N_I,
  TX_CLK_I               => TX_CLK_I,

  TX_POLARITY_I          => TX_POLARITY_I,
  TX_PRBS_SEL_I          => TX_PRBS_SEL_I, -- 3-bit
  TX_PRBS_FORCE_ERR_I    => TX_PRBS_FORCE_ERR_I,
  TX_8B10B_EN_I          => TX_8B10B_EN_I,
  TX_8B10B_BYPASS_I      => TX_8B10B_BYPASS_I, -- 8-bit
  TX_CHAR_IS_K_I         => TX_CHAR_IS_K_I, -- 8-bit
  TX_CHAR_DISPMODE_I     => TX_CHAR_DISPMODE_I, -- 8-bit
  TX_CHAR_DISPVAL_I      => TX_CHAR_DISPVAL_I, -- 8-bit
  TX_ELEC_IDLE_I         => TX_ELEC_IDLE_I,
  TX_DETECT_RX_I         => TX_DETECT_RX_I,

  TX_DATA_I              => TX_DATA_I, -- 64-bit

  TX_RESET_DONE_O        => TX_RESET_DONE_O,
  TX_BUF_ERR_O           => TX_BUF_ERR_O,
  TX_DETECT_RX_PRESENT_O => TX_DETECT_RX_PRESENT_O,
  TX_DETECT_RX_DONE_O    => TX_DETECT_RX_DONE_O,

  -- Receiver
  RX_RESET_I           => RX_RESET_I,
  RX_PMA_RESET_I       => RX_PMA_RESET_I,
  RX_EQA_RESET_I       => RX_EQA_RESET_I,
  RX_CDR_RESET_I       => RX_CDR_RESET_I,
  RX_PCS_RESET_I       => RX_PCS_RESET_I,
  RX_BUF_RESET_I       => RX_BUF_RESET_I,
  RX_POWER_DOWN_N_I    => RX_POWER_DOWN_N_I,
  RX_CLK_I             => RX_CLK_I,

  RX_POLARITY_I        => RX_POLARITY_I,
  RX_PRBS_SEL_I        => RX_PRBS_SEL_I, -- 3-bit
  RX_PRBS_CNT_RESET_I  => RX_PRBS_CNT_RESET_I,
  RX_8B10B_EN_I        => RX_8B10B_EN_I,
  RX_8B10B_BYPASS_I    => RX_8B10B_BYPASS_I, -- 8-bit
  RX_EN_EI_DETECTOR_I  => RX_EN_EI_DETECTOR_I,
  RX_COMMA_DETECT_EN_I => RX_COMMA_DETECT_EN_I,
  RX_SLIDE_I           => RX_SLIDE_I,
  RX_MCOMMA_ALIGN_I    => RX_MCOMMA_ALIGN_I,
  RX_PCOMMA_ALIGN_I    => RX_PCOMMA_ALIGN_I,

  RX_CLK_O             => RX_CLK_O,

  RX_NOT_IN_TABLE_O    => RX_NOT_IN_TABLE_O, -- 8-bit
  RX_CHAR_IS_COMMA_O   => RX_CHAR_IS_COMMA_O, -- 8-bit
  RX_CHAR_IS_K_O       => RX_CHAR_IS_K_O, -- 8-bit
  RX_DISP_ERR_O        => RX_DISP_ERR_O, -- 8-bit
  RX_PRBS_ERR_O        => RX_PRBS_ERR_O,
  RX_BUF_ERR_O         => RX_BUF_ERR_O,
  RX_BYTE_IS_ALIGNED_O => RX_BYTE_IS_ALIGNED_O,
  RX_BYTE_REALIGN_O    => RX_BYTE_REALIGN_O,
  RX_RESET_DONE_O      => RX_RESET_DONE_O,
  RX_EI_EN_O           => RX_EI_EN_O,

  RX_DATA_O            => RX_DATA_O, -- 64-bit

  -- Register File
  REGFILE_CLK_I        => REGFILE_CLK_I,
  REGFILE_WE_I         => REGFILE_WE_I,
  REGFILE_EN_I         => REGFILE_EN_I,
  REGFILE_ADDR_I       => REGFILE_ADDR_I, -- 8-bit
  REGFILE_DI_I         => REGFILE_DI_I, -- 16-bit
  REGFILE_MASK_I       => REGFILE_MASK_I, -- 16-bit

  REGFILE_DO_O         => REGFILE_DO_O, -- 16-bit
  REGFILE_RDY_O        => REGFILE_RDY_O,

  -- ADPLL
  PLL_RESET_I          => PLL_RESET_I,
  PLL_CLK_O            => PLL_CLK_O,

  -- Miscellaneous
  LOOPBACK_I           => LOOPBACK_I, -- 3-bit
);
