//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 May 2024)
//  Compile Time: 1970-01-01 00:59:59
//  Program Run:  2024-07-11 21:35:55
//  Program Call: p_r +sp -i /home/user/FPGA/Boards/GateMate/gatemate_ila/net/ila_top_synth24-07-11_21-35-27.v -o /home/user/FPGA/Boards/GateMate/gatemate_ila/p_r_out/ila_top_24-07-11_21-35-27 -sp -cCP +uCIO -ccf /home/user/FPGA/Boards/GateMate/gatemate_ila/src/ILA_top.ccf 
//  File Type:    Verilog

// Gatecount:    277
module ila_top_24-07-11_21-35-27 (clk , i_mosi_ILA , i_sclk_ILA , i_ss_ILA ,
       led , o_miso_ILA 
       ) ;

input  clk;
input  i_mosi_ILA;
input  i_sclk_ILA;
input  i_ss_ILA;

output led;
output o_miso_ILA;



wire clk;
wire led;
wire na1_1;
wire na1_1_i;
wire na1_2;
wire na1_2_i;
wire na2_1;
wire na2_1_i;
wire na2_2;
wire na2_2_i;
wire na3_1;
wire na3_1_i;
wire na3_2;
wire na3_2_i;
wire na4_1;
wire na4_1_i;
wire na4_2;
wire na4_2_i;
wire na5_1;
wire na5_1_i;
wire na6_2;
wire na6_2_i;
wire na7_1;
wire na8_1;
wire na9_1;
wire na9_1_i;
wire na10_1;
wire na10_1_i;
wire na10_2;
wire na10_2_i;
wire na11_1;
wire na11_1_i;
wire na13_2;
wire na13_2_i;
wire na14_1;
wire na14_1_i;
wire na14_2;
wire na14_2_i;
wire na16_1;
wire na16_1_i;
wire na16_2;
wire na16_2_i;
wire na17_1;
wire na17_1_i;
wire na17_2;
wire na17_2_i;
wire na18_1;
wire na18_1_i;
wire na18_2;
wire na18_2_i;
wire na19_2;
wire na19_2_i;
wire na20_2;
wire na21_1;
wire na21_1_i;
wire na23_1;
wire na23_1_i;
wire na23_2;
wire na23_2_i;
wire na25_1;
wire na25_1_i;
wire na25_2;
wire na25_2_i;
wire na27_1;
wire na27_1_i;
wire na27_2;
wire na27_2_i;
wire na28_1;
wire na28_1_i;
wire na28_2;
wire na28_2_i;
wire na29_1;
wire na29_1_i;
wire na29_2;
wire na29_2_i;
wire na33_1;
wire na33_1_i;
wire na33_2;
wire na33_2_i;
wire na34_1;
wire na34_1_i;
wire na34_2;
wire na34_2_i;
wire na35_1;
wire na35_1_i;
wire na36_1;
wire na36_1_i;
wire na36_2;
wire na36_2_i;
wire na37_1;
wire na37_1_i;
wire na37_2;
wire na37_2_i;
wire na39_2;
wire na39_2_i;
wire na40_1;
wire na40_1_i;
wire na41_1;
wire na41_1_i;
wire na41_2;
wire na41_2_i;
wire na43_1;
wire na43_1_i;
wire na44_1;
wire na44_1_i;
wire na44_2;
wire na44_2_i;
wire na45_1;
wire na45_1_i;
wire na47_1;
wire na47_1_i;
wire na47_2;
wire na47_2_i;
wire na48_1;
wire na48_1_i;
wire na49_2;
wire na51_1;
wire na51_1_i;
wire na51_2;
wire na51_2_i;
wire na52_1;
wire na52_1_i;
wire na52_2;
wire na52_2_i;
wire na53_1;
wire na53_1_i;
wire na54_2;
wire na54_2_i;
wire na55_1;
wire na56_1;
wire na56_1_i;
wire na57_1;
wire na57_1_i;
wire na58_1;
wire na58_1_i;
wire na58_2;
wire na58_2_i;
wire na59_1;
wire na59_1_i;
wire na59_2;
wire na59_2_i;
wire na61_1;
wire na61_1_i;
wire na61_2;
wire na61_2_i;
wire na63_1;
wire na63_1_i;
wire na65_1;
wire na65_1_i;
wire na66_1;
wire na66_1_i;
wire na66_2;
wire na66_2_i;
wire na67_1;
wire na67_1_i;
wire na68_1;
wire na68_1_i;
wire na69_1;
wire na69_1_i;
wire na75_1;
wire na75_1_i;
wire na79_1;
wire na79_1_i;
wire na80_1;
wire na80_1_i;
wire na81_1;
wire na81_1_i;
wire na82_1;
wire na82_1_i;
wire na83_1;
wire na83_1_i;
wire na84_1;
wire na84_1_i;
wire na85_1;
wire na85_1_i;
wire na86_1;
wire na86_1_i;
wire na87_1;
wire na87_1_i;
wire na88_1;
wire na88_1_i;
wire na89_1;
wire na89_1_i;
wire na90_1;
wire na90_1_i;
wire na90_2;
wire na90_2_i;
wire na93_1;
wire na93_1_i;
wire na93_2;
wire na93_2_i;
wire na94_1;
wire na94_1_i;
wire na94_2;
wire na94_2_i;
wire na97_2;
wire na97_2_i;
wire na99_1;
wire na99_1_i;
wire na100_2;
wire na100_2_i;
wire na101_1;
wire na101_1_i;
wire na101_2;
wire na101_2_i;
wire na103_1;
wire na103_1_i;
wire na103_2;
wire na103_2_i;
wire na105_1;
wire na105_1_i;
wire na106_2;
wire na106_2_i;
wire na107_1;
wire na107_1_i;
wire na112_2;
wire na112_2_i;
wire na113_2;
wire na114_1;
wire na115_1;
wire na115_1_i;
wire na115_2;
wire na115_2_i;
wire na116_2;
wire na116_2_i;
wire na117_1;
wire na121_1;
wire na122_1;
wire na122_1_i;
wire na123_1;
wire na124_1;
wire na124_1_i;
wire na125_1;
wire na126_1;
wire na126_1_i;
wire na129_1;
wire na129_2;
wire na129_4;
wire na131_1;
wire na131_2;
wire na131_4;
wire na133_1;
wire na133_2;
wire na133_4;
wire na135_1;
wire na135_2;
wire na135_4;
wire na137_1;
wire na137_2;
wire na137_4;
wire na138_1;
wire na138_2;
wire na138_4;
wire na140_1;
wire na140_2;
wire na140_4;
wire na142_1;
wire na142_2;
wire na145_1;
wire na145_2;
wire na145_4;
wire na147_1;
wire na147_2;
wire na147_4;
wire na149_1;
wire na149_2;
wire na149_4;
wire na151_1;
wire na151_2;
wire na151_4;
wire na152_1;
wire na152_4;
wire na153_1;
wire na153_2;
wire na153_4;
wire na155_1;
wire na155_2;
wire na155_4;
wire na157_1;
wire na157_2;
wire na157_4;
wire na159_1;
wire na159_2;
wire na159_4;
wire na161_1;
wire na162_1;
wire na162_4;
wire na163_1;
wire na163_2;
wire na163_4;
wire na165_1;
wire na165_2;
wire na165_4;
wire na167_1;
wire na167_2;
wire na167_4;
wire na169_1;
wire na169_2;
wire na169_4;
wire na171_1;
wire na172_1;
wire na172_4;
wire na173_1;
wire na173_2;
wire na173_4;
wire na175_1;
wire na175_2;
wire na175_4;
wire na177_1;
wire na177_2;
wire na177_4;
wire na179_1;
wire na179_2;
wire na179_4;
wire na181_1;
wire na182_1;
wire na182_4;
wire na183_1;
wire na183_2;
wire na183_4;
wire na185_1;
wire na185_2;
wire na185_4;
wire na187_1;
wire na187_2;
wire na187_4;
wire na189_1;
wire na189_2;
wire na189_4;
wire na191_1;
wire na194_1;
wire na194_2;
wire na211_1;
wire na211_1_i;
wire na212_2;
wire na212_2_i;
wire na262_1;
wire na262_1_i;
wire na273_2;
wire na273_2_i;
wire na309_1;
wire na310_1;
wire na311_1;
wire na312_1;
wire na315_3;
wire na315_4;
wire na315_5;
wire na315_6;
wire na316_3;
wire na316_4;
wire na316_5;
wire na316_6;
wire na318_1;
wire na319_1;
wire na320_1;
wire na321_1;
wire na322_1;
wire na322_2;
wire na323_2;
wire na324_1;
wire na325_1;
wire na325_9;
wire na326_1;
wire na327_1;
wire na328_1;
wire na329_1;
wire na330_1;
wire na331_2;
wire na332_1;
wire na333_1;
wire na334_1;
wire na335_1;
wire na336_2;
wire na337_1;
wire na338_1;
wire na339_1;
wire na340_1;
wire na341_2;
wire na342_1;
wire na343_1;
wire na343_9;
wire na344_1;
wire na345_1;
wire na346_2;
wire na347_1;
wire na348_1;
wire na349_1;
wire na349_9;
wire na350_2;
wire na351_1;
wire na352_1;
wire na353_1;
wire na354_1;
wire na355_1;
wire na356_1;
wire na357_1;
wire na358_1;
wire na359_1;
wire na360_1;
wire na360_9;
wire na361_2;
wire na362_1;
wire na363_1;
wire na363_9;
wire na364_1;
wire na365_2;
wire na366_1;
wire na367_1;
wire na368_1;
wire na369_1;
wire na369_9;
wire na370_1;
wire na371_1;
wire na371_4;
wire na372_2;
wire na373_2;
wire na374_2;
wire na375_1;
wire na375_9;
wire na376_2;
wire na377_1;
wire na377_9;
wire na378_2;
wire na379_1;
wire na379_9;
wire na380_2;
wire na381_1;
wire na381_9;
wire na382_2;
wire na383_1;
wire na383_9;
wire na384_2;
wire na385_1;
wire na385_9;
wire na386_2;
wire na387_1;
wire na387_9;
wire na388_2;
wire na389_1;
wire na389_9;
wire na390_2;
wire na391_1;
wire na391_9;
wire na392_2;
wire na393_1;
wire na393_9;
wire na394_2;
wire na395_1;
wire na395_9;
wire na396_2;
wire na397_1;
wire na397_9;
wire na398_2;
wire na399_1;
wire na399_9;
wire na400_2;
wire na401_1;
wire na401_9;
wire na402_2;
wire na403_1;
wire na403_9;
wire na404_2;
wire na405_1;
wire na405_9;
wire na406_2;
wire na407_1;
wire na407_9;
wire na408_2;
wire na409_1;
wire na409_9;
wire na410_2;
wire na411_1;
wire na411_9;
wire na412_2;
wire na413_1;
wire na413_9;
wire na414_2;
wire na415_1;
wire na415_9;
wire na416_2;
wire na417_1;
wire na417_9;
wire na418_2;
wire na419_1;
wire na419_9;
wire na420_2;
wire na421_1;
wire na421_9;
wire na422_2;
wire na423_1;
wire na423_9;
wire na424_2;
wire na425_1;
wire na425_9;
wire na426_2;
wire na427_1;
wire na427_9;
wire na428_2;
wire na429_1;
wire na429_9;
wire na430_2;
wire na431_1;
wire na432_2;
wire na433_2;
wire na434_2;
wire na435_2;
wire na436_2;
wire na437_2;
wire na438_2;
wire na439_2;
wire na440_2;
wire na441_2;
wire na442_2;
wire na443_2;
wire na444_2;
wire na445_2;
wire na446_2;
wire na447_2;
wire na448_2;
wire na449_2;
wire na450_2;
wire na451_2;
wire na452_2;
wire na453_2;
wire na454_2;
wire na455_2;
wire na456_2;
wire na457_2;
wire na458_2;
wire na459_2;
wire na460_2;
wire na461_2;
wire i_ss_ILA;
wire na331_10;
wire na336_10;
wire na346_10;
wire na350_10;
wire na361_10;
wire na365_10;
wire na372_10;
wire na373_10;
wire na374_10;
wire na376_10;
wire na378_10;
wire na380_10;
wire na382_10;
wire na384_10;
wire na386_10;
wire na388_10;
wire na390_10;
wire na392_10;
wire na394_10;
wire na396_10;
wire na398_10;
wire na400_10;
wire na402_10;
wire na404_10;
wire na406_10;
wire na408_10;
wire na410_10;
wire na412_10;
wire na414_10;
wire na416_10;
wire na418_10;
wire na420_10;
wire na422_10;
wire na424_10;
wire na426_10;
wire na428_10;
wire na430_10;
wire na317_120;
wire i_mosi_ILA;
wire i_sclk_ILA;
wire o_miso_ILA;

// C_AND/D//AND/D      x35y53     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1_1 ( .OUT(na1_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(na129_2), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1_2 ( .OUT(na1_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1_4 ( .OUT(na1_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(na129_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1_5 ( .OUT(na1_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1_2_i) );
// C_AND/D//ORAND/D      x39y39     80'h00_FE00_80_0000_0C88_AACE
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2_1 ( .OUT(na2_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2_2), .IN6(1'b1), .IN7(na431_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2_2 ( .OUT(na2_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a2_4 ( .OUT(na2_2_i), .IN1(na2_2), .IN2(na364_1), .IN3(1'b0), .IN4(na21_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2_5 ( .OUT(na2_2), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2_2_i) );
// C_AND/D//AND/D      x46y48     80'h00_FE00_80_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3_1 ( .OUT(na3_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(na319_1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3_2 ( .OUT(na3_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3_4 ( .OUT(na3_2_i), .IN1(na324_1), .IN2(1'b1), .IN3(1'b1), .IN4(na452_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3_5 ( .OUT(na3_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3_2_i) );
// C_AND/D//AND/D      x40y47     80'h00_FE00_80_0000_0C88_58CF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4_1 ( .OUT(na4_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na67_1), .IN6(na75_1), .IN7(~na4_2), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4_2 ( .OUT(na4_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4_4 ( .OUT(na4_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na94_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4_5 ( .OUT(na4_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4_2_i) );
// C_AND/D///      x36y35     80'h00_FD00_00_0000_0C88_34FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5_1 ( .OUT(na5_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na8_1), .IN6(na7_1), .IN7(1'b1), .IN8(~na312_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5_2 ( .OUT(na5_1), .CLK(~na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5_1_i) );
// C_///AND/D      x39y40     80'h00_FD00_80_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6_4 ( .OUT(na6_2_i), .IN1(1'b1), .IN2(na7_1), .IN3(1'b1), .IN4(~na312_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6_5 ( .OUT(na6_2), .CLK(~na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6_2_i) );
// C_AND////      x39y36     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7_1 ( .OUT(na7_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na448_2), .IN6(na66_2), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x39y41     80'h00_0018_00_0040_0C33_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1), .IN1(~na320_1), .IN2(~na10_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na51_2), .IN7(1'b0), .IN8(1'b0),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x39y42     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9_1 ( .OUT(na9_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(1'b1), .IN7(na321_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a9_2 ( .OUT(na9_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na9_1_i) );
// C_AND/D//AND/D      x41y42     80'h00_FE00_80_0000_0C88_3C3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a10_1 ( .OUT(na10_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na310_1), .IN7(1'b1), .IN8(~na312_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a10_2 ( .OUT(na10_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na10_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a10_4 ( .OUT(na10_2_i), .IN1(1'b1), .IN2(na10_1), .IN3(1'b1), .IN4(~na312_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a10_5 ( .OUT(na10_2), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na10_2_i) );
// C_AND/D///      x38y38     80'h00_FE00_00_0000_0888_3C42
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a11_1 ( .OUT(na11_1_i), .IN1(na40_1), .IN2(~na63_1), .IN3(~na45_1), .IN4(na65_1), .IN5(1'b1), .IN6(na6_2), .IN7(1'b1), .IN8(~na68_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a11_2 ( .OUT(na11_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na11_1_i) );
// C_///AND/D      x39y48     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a13_4 ( .OUT(na13_2_i), .IN1(na67_1), .IN2(1'b1), .IN3(na4_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a13_5 ( .OUT(na13_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na13_2_i) );
// C_AND/D//AND/D      x39y56     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a14_1 ( .OUT(na14_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(na142_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a14_2 ( .OUT(na14_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na14_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a14_4 ( .OUT(na14_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(na142_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a14_5 ( .OUT(na14_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na14_2_i) );
// C_AND/D//AND/D      x35y49     80'h00_FE00_80_0000_0C88_A2F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a16_1 ( .OUT(na16_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na67_1), .IN6(~na75_1), .IN7(na4_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a16_2 ( .OUT(na16_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na16_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a16_4 ( .OUT(na16_2_i), .IN1(na67_1), .IN2(na435_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a16_5 ( .OUT(na16_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na16_2_i) );
// C_AND/D//AND/D      x41y41     80'h00_FE00_80_0000_0C88_3C3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a17_1 ( .OUT(na17_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na10_2), .IN7(1'b1), .IN8(~na312_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a17_2 ( .OUT(na17_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na17_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a17_4 ( .OUT(na17_2_i), .IN1(na17_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na312_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a17_5 ( .OUT(na17_2), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na17_2_i) );
// C_AND/D//AND/D      x42y44     80'h00_FE00_80_0000_0C88_38CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a18_1 ( .OUT(na18_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(na273_2), .IN7(1'b1), .IN8(~na18_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a18_2 ( .OUT(na18_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na18_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a18_4 ( .OUT(na18_2_i), .IN1(na328_1), .IN2(1'b1), .IN3(1'b1), .IN4(na452_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a18_5 ( .OUT(na18_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na18_2_i) );
// C_///ICOMP/D      x39y45     80'h00_FE00_80_0000_0C08_FFC6
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a19_4 ( .OUT(na19_2_i), .IN1(na19_2), .IN2(~na20_2), .IN3(1'b0), .IN4(~na21_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a19_5 ( .OUT(na19_2), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na19_2_i) );
// C_///AND/      x39y42     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a20_4 ( .OUT(na20_2), .IN1(1'b1), .IN2(na6_2), .IN3(na45_1), .IN4(na57_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x36y46     80'h00_FE00_00_0000_0888_EF5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a21_1 ( .OUT(na21_1_i), .IN1(1'b0), .IN2(na323_2), .IN3(~na69_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na211_1), .IN8(na21_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a21_2 ( .OUT(na21_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na21_1_i) );
// C_AND/D//AND/D      x36y50     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a23_1 ( .OUT(na23_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(na145_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a23_2 ( .OUT(na23_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na23_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a23_4 ( .OUT(na23_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(na145_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a23_5 ( .OUT(na23_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na23_2_i) );
// C_ORAND/D//AND/D      x43y46     80'h00_FE00_80_0000_0C88_EA82
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a25_1 ( .OUT(na25_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(1'b0), .IN7(na439_2), .IN8(na18_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a25_2 ( .OUT(na25_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na25_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a25_4 ( .OUT(na25_2_i), .IN1(na106_2), .IN2(~na51_2), .IN3(na112_2), .IN4(na440_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a25_5 ( .OUT(na25_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na25_2_i) );
// C_AND/D//AND/D      x41y45     80'h00_FE00_80_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na326_1), .IN6(1'b1), .IN7(1'b1), .IN8(na452_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a27_2 ( .OUT(na27_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na27_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a27_4 ( .OUT(na27_2_i), .IN1(na106_2), .IN2(na327_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a27_5 ( .OUT(na27_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na27_2_i) );
// C_AND/D//AND/D      x37y53     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a28_1 ( .OUT(na28_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(1'b1), .IN8(na135_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a28_2 ( .OUT(na28_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na28_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a28_4 ( .OUT(na28_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(1'b1), .IN4(na135_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a28_5 ( .OUT(na28_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na28_2_i) );
// C_AND/D//AND/D      x37y55     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a29_1 ( .OUT(na29_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(1'b1), .IN8(na140_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a29_2 ( .OUT(na29_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na29_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a29_4 ( .OUT(na29_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(1'b1), .IN4(na140_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a29_5 ( .OUT(na29_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na29_2_i) );
// C_AND/D//AND/D      x39y55     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_1 ( .OUT(na33_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(na137_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a33_2 ( .OUT(na33_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na33_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a33_4 ( .OUT(na33_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(na137_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a33_5 ( .OUT(na33_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na33_2_i) );
// C_AND/D//AND/D      x42y45     80'h00_FE00_80_0000_0C88_4AAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a34_1 ( .OUT(na34_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na262_1), .IN6(1'b1), .IN7(~na34_2), .IN8(na452_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a34_2 ( .OUT(na34_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na34_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a34_4 ( .OUT(na34_2_i), .IN1(na106_2), .IN2(1'b1), .IN3(na352_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a34_5 ( .OUT(na34_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na34_2_i) );
// C_AND/D///      x34y44     80'h00_FE00_00_0000_0888_3C44
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a35_1 ( .OUT(na35_1_i), .IN1(~na40_1), .IN2(na63_1), .IN3(~na45_1), .IN4(na65_1), .IN5(1'b1), .IN6(na6_2), .IN7(1'b1), .IN8(~na68_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a35_2 ( .OUT(na35_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na35_1_i) );
// C_AND/D//AND/D      x39y53     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(na133_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a36_2 ( .OUT(na36_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na36_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a36_4 ( .OUT(na36_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(na133_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a36_5 ( .OUT(na36_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na36_2_i) );
// C_AND/D//AND/D      x37y51     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a37_1 ( .OUT(na37_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(na149_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a37_2 ( .OUT(na37_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na37_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a37_4 ( .OUT(na37_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(na149_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a37_5 ( .OUT(na37_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na37_2_i) );
// C_///AND/D      x37y50     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a39_4 ( .OUT(na39_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(1'b1), .IN4(na138_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a39_5 ( .OUT(na39_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na39_2_i) );
// C_MX4b/D///      x41y43     80'h00_FD00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a40_1 ( .OUT(na40_1_i), .IN1(1'b1), .IN2(na7_1), .IN3(1'b1), .IN4(na312_1), .IN5(na40_1), .IN6(na10_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a40_2 ( .OUT(na40_1), .CLK(~na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na40_1_i) );
// C_AND/D//AND/D      x40y53     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a41_1 ( .OUT(na41_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(1'b1), .IN8(na151_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a41_2 ( .OUT(na41_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na41_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a41_4 ( .OUT(na41_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(1'b1), .IN4(na151_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a41_5 ( .OUT(na41_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na41_2_i) );
// C_AND/D///      x43y44     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a43_1 ( .OUT(na43_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(1'b1), .IN7(na329_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a43_2 ( .OUT(na43_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na43_1_i) );
// C_AND/D//AND/D      x43y43     80'h00_FE00_80_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a44_1 ( .OUT(na44_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(na330_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a44_2 ( .OUT(na44_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na44_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a44_4 ( .OUT(na44_2_i), .IN1(na106_2), .IN2(1'b1), .IN3(1'b1), .IN4(na332_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a44_5 ( .OUT(na44_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na44_2_i) );
// C_ORAND/D///      x38y39     80'h00_FE00_00_0000_0888_EFC5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1_i), .IN1(~na106_2), .IN2(1'b0), .IN3(1'b0), .IN4(na21_1), .IN5(1'b1), .IN6(1'b1), .IN7(na45_1), .IN8(na11_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_2 ( .OUT(na45_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na45_1_i) );
// C_AND/D//AND/D      x43y42     80'h00_FE00_80_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a47_1 ( .OUT(na47_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(1'b1), .IN7(1'b1), .IN8(na333_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a47_2 ( .OUT(na47_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na47_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a47_4 ( .OUT(na47_2_i), .IN1(na106_2), .IN2(1'b1), .IN3(1'b1), .IN4(na335_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a47_5 ( .OUT(na47_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na47_2_i) );
// C_AND/D///      x36y43     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a48_1 ( .OUT(na48_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na438_2), .IN6(1'b1), .IN7(1'b1), .IN8(na334_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a48_2 ( .OUT(na48_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na48_1_i) );
// C_///AND/      x37y44     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a49_4 ( .OUT(na49_2), .IN1(na19_2), .IN2(na6_2), .IN3(na45_1), .IN4(na57_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP/D//ORAND/D      x39y44     80'h00_FE00_80_0000_0C88_9AEA
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a51_1 ( .OUT(na51_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na106_2), .IN6(1'b0), .IN7(~na445_2), .IN8(~na444_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a51_2 ( .OUT(na51_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na51_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a51_4 ( .OUT(na51_2_i), .IN1(na106_2), .IN2(1'b0), .IN3(na34_1), .IN4(na446_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a51_5 ( .OUT(na51_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na51_2_i) );
// C_AND/D//AND/D      x42y47     80'h00_FE00_80_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a52_1 ( .OUT(na52_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na337_1), .IN6(1'b1), .IN7(1'b1), .IN8(na452_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a52_2 ( .OUT(na52_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na52_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a52_4 ( .OUT(na52_2_i), .IN1(na106_2), .IN2(na362_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a52_5 ( .OUT(na52_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na52_2_i) );
// C_AND/D///      x36y44     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a53_1 ( .OUT(na53_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(na338_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a53_2 ( .OUT(na53_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na53_1_i) );
// C_///AND/D      x37y47     80'h00_FE00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a54_4 ( .OUT(na54_2_i), .IN1(na339_1), .IN2(1'b1), .IN3(1'b1), .IN4(na21_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a54_5 ( .OUT(na54_2), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na54_2_i) );
// C_AND////      x39y43     80'h00_0018_00_0000_0C88_28FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na19_2), .IN6(na6_2), .IN7(na45_1), .IN8(~na57_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x40y43     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a56_1 ( .OUT(na56_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na340_1), .IN6(1'b1), .IN7(1'b1), .IN8(na21_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a56_2 ( .OUT(na56_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na56_1_i) );
// C_MX4a/D///      x36y40     80'h00_FE00_00_0040_0C0C_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a57_1 ( .OUT(na57_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na341_2), .IN4(na57_1), .IN5(1'b1), .IN6(~na442_2), .IN7(1'b1), .IN8(na21_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a57_2 ( .OUT(na57_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na57_1_i) );
// C_AND/D//AND/D      x34y41     80'h00_FE00_80_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a58_1 ( .OUT(na58_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(na342_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a58_2 ( .OUT(na58_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na58_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a58_4 ( .OUT(na58_2_i), .IN1(na106_2), .IN2(1'b1), .IN3(na344_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a58_5 ( .OUT(na58_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na58_2_i) );
// C_AND/D//AND/D      x36y52     80'h00_FE00_80_0000_0C88_CC3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a59_1 ( .OUT(na59_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(1'b1), .IN8(na138_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a59_2 ( .OUT(na59_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na59_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a59_4 ( .OUT(na59_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(1'b1), .IN4(~na59_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a59_5 ( .OUT(na59_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na59_2_i) );
// C_AND/D//AND/D      x37y49     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a61_1 ( .OUT(na61_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(1'b1), .IN8(na147_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a61_2 ( .OUT(na61_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na61_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a61_4 ( .OUT(na61_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(1'b1), .IN4(na147_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a61_5 ( .OUT(na61_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na61_2_i) );
// C_MX4b/D///      x41y40     80'h00_FD00_00_0040_0A30_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a63_1 ( .OUT(na63_1_i), .IN1(1'b1), .IN2(~na7_1), .IN3(1'b1), .IN4(na312_1), .IN5(na17_1), .IN6(na63_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a63_2 ( .OUT(na63_1), .CLK(~na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na63_1_i) );
// C_MX4b/D///      x44y38     80'h00_FD00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a65_1 ( .OUT(na65_1_i), .IN1(1'b1), .IN2(~na7_1), .IN3(1'b1), .IN4(~na312_1), .IN5(1'b0), .IN6(1'b0), .IN7(na436_2), .IN8(na65_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a65_2 ( .OUT(na65_1), .CLK(~na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na65_1_i) );
// C_AND*/D//ICOMP*/D      x39y34     80'h00_FE00_80_0000_0387_3C39
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a66_1 ( .OUT(na66_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na66_1), .IN7(1'b1), .IN8(~na312_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a66_2 ( .OUT(na66_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na66_1_i) );
C_ICOMP    #(.CPE_CFG (9'b1_1000_0000)) 
           _a66_4 ( .OUT(na66_2_i), .IN1(~na449_2), .IN2(~na66_1), .IN3(1'b0), .IN4(na312_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a66_5 ( .OUT(na66_2), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na66_2_i) );
// C_ORAND/D///      x35y47     80'h00_FE00_00_0000_0888_FE5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_1 ( .OUT(na67_1_i), .IN1(1'b0), .IN2(na323_2), .IN3(~na69_1), .IN4(1'b0), .IN5(na67_1), .IN6(na212_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a67_2 ( .OUT(na67_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na67_1_i) );
// C_MX4b/D///      x34y38     80'h00_FD00_00_0040_0AC0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a68_1 ( .OUT(na68_1_i), .IN1(1'b1), .IN2(~na7_1), .IN3(1'b1), .IN4(~na312_1), .IN5(1'b0), .IN6(1'b0), .IN7(na434_2), .IN8(na68_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a68_2 ( .OUT(na68_1), .CLK(~na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na68_1_i) );
// C_AND/D///      x36y41     80'h00_FE00_00_0000_0888_CC14
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a69_1 ( .OUT(na69_1_i), .IN1(~na40_1), .IN2(na63_1), .IN3(~na45_1), .IN4(~na65_1), .IN5(1'b1), .IN6(na6_2), .IN7(1'b1),
                    .IN8(na68_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a69_2 ( .OUT(na69_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na69_1_i) );
// C_MX2b/D///      x39y50     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1_i), .IN1(~na67_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4_2), .IN8(na94_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a75_2 ( .OUT(na75_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na75_1_i) );
// C_MX2b/D///      x42y35     80'h00_F600_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a79_1 ( .OUT(na79_1_i), .IN1(1'b1), .IN2(~na6_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na79_1), .IN8(~na115_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a79_2 ( .OUT(na79_1), .CLK(na311_1), .EN(~na117_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na79_1_i) );
// C_MX2b/D///      x43y36     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1_i), .IN1(1'b1), .IN2(~na6_2), .IN3(1'b0), .IN4(1'b0), .IN5(na153_1), .IN6(na453_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a80_2 ( .OUT(na80_1), .CLK(na311_1), .EN(~na117_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na80_1_i) );
// C_MX2b/D///      x41y36     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a81_1 ( .OUT(na81_1_i), .IN1(1'b1), .IN2(~na6_2), .IN3(1'b0), .IN4(1'b0), .IN5(na153_2), .IN6(na454_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a81_2 ( .OUT(na81_1), .CLK(na311_1), .EN(~na117_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na81_1_i) );
// C_MX2b/D///      x42y38     80'h00_F600_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a82_1 ( .OUT(na82_1_i), .IN1(1'b1), .IN2(na6_2), .IN3(1'b0), .IN4(1'b0), .IN5(na455_2), .IN6(na155_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a82_2 ( .OUT(na82_1), .CLK(na311_1), .EN(~na117_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na82_1_i) );
// C_MX2b/D///      x42y39     80'h00_F600_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a83_1 ( .OUT(na83_1_i), .IN1(1'b1), .IN2(na6_2), .IN3(1'b0), .IN4(1'b0), .IN5(na456_2), .IN6(na155_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a83_2 ( .OUT(na83_1), .CLK(na311_1), .EN(~na117_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na83_1_i) );
// C_MX2b/D///      x43y39     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a84_1 ( .OUT(na84_1_i), .IN1(1'b1), .IN2(~na6_2), .IN3(1'b0), .IN4(1'b0), .IN5(na157_1), .IN6(na457_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a84_2 ( .OUT(na84_1), .CLK(na311_1), .EN(~na117_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na84_1_i) );
// C_MX2b/D///      x43y37     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a85_1 ( .OUT(na85_1_i), .IN1(1'b1), .IN2(~na6_2), .IN3(1'b0), .IN4(1'b0), .IN5(na157_2), .IN6(na458_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a85_2 ( .OUT(na85_1), .CLK(na311_1), .EN(~na117_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na85_1_i) );
// C_MX2b/D///      x43y41     80'h00_F600_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a86_1 ( .OUT(na86_1_i), .IN1(1'b1), .IN2(na6_2), .IN3(1'b0), .IN4(1'b0), .IN5(na459_2), .IN6(na159_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a86_2 ( .OUT(na86_1), .CLK(na311_1), .EN(~na117_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na86_1_i) );
// C_MX2b/D///      x39y38     80'h00_F600_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a87_1 ( .OUT(na87_1_i), .IN1(1'b1), .IN2(na6_2), .IN3(1'b0), .IN4(1'b0), .IN5(na460_2), .IN6(na159_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a87_2 ( .OUT(na87_1), .CLK(na311_1), .EN(~na117_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na87_1_i) );
// C_MX2b/D///      x44y39     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a88_1 ( .OUT(na88_1_i), .IN1(1'b1), .IN2(~na6_2), .IN3(1'b0), .IN4(1'b0), .IN5(na161_1), .IN6(na461_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a88_2 ( .OUT(na88_1), .CLK(na311_1), .EN(~na117_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na88_1_i) );
// C_ICOMP/D///      x42y50     80'h00_FE00_00_0000_0C88_6AFF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na106_2), .IN6(1'b0), .IN7(~na441_2), .IN8(na89_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a89_2 ( .OUT(na89_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_1_i) );
// C_AND/D//AND/D      x35y41     80'h00_FE00_80_0000_0C88_CAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(1'b1), .IN7(1'b1), .IN8(na347_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a90_2 ( .OUT(na90_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na90_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a90_4 ( .OUT(na90_2_i), .IN1(na106_2), .IN2(1'b1), .IN3(na348_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a90_5 ( .OUT(na90_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na90_2_i) );
// C_AND/D//AND/D      x40y54     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_1 ( .OUT(na93_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na323_2), .IN7(1'b1), .IN8(na131_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a93_2 ( .OUT(na93_1), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na93_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a93_4 ( .OUT(na93_2_i), .IN1(1'b1), .IN2(na323_2), .IN3(1'b1), .IN4(na131_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a93_5 ( .OUT(na93_2), .CLK(na194_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na93_2_i) );
// C_AND/D//AND/D      x40y48     80'h00_FE00_80_0000_0C88_41AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a94_1 ( .OUT(na94_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na54_2), .IN6(~na97_2), .IN7(~na56_1), .IN8(na94_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a94_2 ( .OUT(na94_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na94_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a94_4 ( .OUT(na94_2_i), .IN1(na309_1), .IN2(1'b1), .IN3(na450_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a94_5 ( .OUT(na94_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na94_2_i) );
// C_///AND/D      x33y44     80'h00_FE00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a97_4 ( .OUT(na97_2_i), .IN1(na438_2), .IN2(1'b1), .IN3(1'b1), .IN4(na351_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a97_5 ( .OUT(na97_2), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na97_2_i) );
// C_AND/D///      x42y48     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a99_1 ( .OUT(na99_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na353_1), .IN6(1'b1), .IN7(1'b1), .IN8(na452_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a99_2 ( .OUT(na99_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na99_1_i) );
// C_///OR/D      x42y48     80'h00_FE00_80_0000_0C0E_FFA5
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a100_4 ( .OUT(na100_2_i), .IN1(~na106_2), .IN2(1'b0), .IN3(na354_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a100_5 ( .OUT(na100_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na100_2_i) );
// C_AND/D//AND/D      x42y49     80'h00_FE00_80_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a101_1 ( .OUT(na101_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(na355_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a101_2 ( .OUT(na101_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na101_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a101_4 ( .OUT(na101_2_i), .IN1(na106_2), .IN2(1'b1), .IN3(1'b1), .IN4(na356_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a101_5 ( .OUT(na101_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na101_2_i) );
// C_AND/D//AND/D      x38y37     80'h00_FE00_80_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_1 ( .OUT(na103_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(na357_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a103_2 ( .OUT(na103_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na103_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a103_4 ( .OUT(na103_2_i), .IN1(na106_2), .IN2(1'b1), .IN3(na358_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a103_5 ( .OUT(na103_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na103_2_i) );
// C_AND/D///      x35y44     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a105_1 ( .OUT(na105_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na359_1), .IN8(na21_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a105_2 ( .OUT(na105_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na105_1_i) );
// C_///ORAND/D      x43y45     80'h00_FE00_80_0000_0C08_FFCE
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a106_4 ( .OUT(na106_2_i), .IN1(na106_2), .IN2(na49_2), .IN3(1'b0), .IN4(na21_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a106_5 ( .OUT(na106_2), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na106_2_i) );
// C_ORAND/D///      x34y39     80'h00_FE00_00_0000_0888_EFC5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a107_1 ( .OUT(na107_1_i), .IN1(~na2_2), .IN2(1'b0), .IN3(1'b0), .IN4(na21_1), .IN5(1'b1), .IN6(1'b1), .IN7(na107_1), .IN8(na35_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a107_2 ( .OUT(na107_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na107_1_i) );
// C_///ORAND/D      x40y45     80'h00_FE00_80_0000_0C08_FFEA
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a112_4 ( .OUT(na112_2_i), .IN1(na67_1), .IN2(1'b0), .IN3(na112_2), .IN4(na113_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a112_5 ( .OUT(na112_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na112_2_i) );
// C_///AND/      x40y46     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a113_4 ( .OUT(na113_2), .IN1(na106_2), .IN2(1'b1), .IN3(1'b1), .IN4(na366_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y45     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a114_1 ( .OUT(na114_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na105_1), .IN7(~na48_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x38y36     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a115_1 ( .OUT(na115_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(1'b1), .IN7(na367_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a115_2 ( .OUT(na115_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na115_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a115_4 ( .OUT(na115_2_i), .IN1(na106_2), .IN2(1'b1), .IN3(na345_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a115_5 ( .OUT(na115_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na115_2_i) );
// C_///AND/D      x33y46     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a116_4 ( .OUT(na116_2_i), .IN1(na106_2), .IN2(na368_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a116_5 ( .OUT(na116_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na116_2_i) );
// C_ORAND////      x46y38     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a117_1 ( .OUT(na117_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2_2), .IN6(~na51_2), .IN7(1'b0), .IN8(~na433_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x38y40     80'h00_0018_00_0040_0A32_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a121_1 ( .OUT(na121_1), .IN1(1'b1), .IN2(~na51_2), .IN3(1'b0), .IN4(1'b0), .IN5(na2_2), .IN6(~na10_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x39y37     80'h00_FD00_00_0040_0AC8_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a122_1 ( .OUT(na122_1_i), .IN1(1'b1), .IN2(na7_1), .IN3(1'b1), .IN4(~na312_1), .IN5(1'b0), .IN6(1'b0), .IN7(na5_1), .IN8(~na121_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a122_2 ( .OUT(na122_1), .CLK(~na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na122_1_i) );
// C_MX2b////      x35y36     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a123_1 ( .OUT(na123_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na446_2), .IN5(na17_1), .IN6(1'b0), .IN7(na370_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x33y36     80'h00_FD00_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a124_1 ( .OUT(na124_1_i), .IN1(1'b1), .IN2(na7_1), .IN3(1'b1), .IN4(na312_1), .IN5(na122_1), .IN6(na123_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a124_2 ( .OUT(na124_1), .CLK(~na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na124_1_i) );
// C_MX2b////      x39y35     80'h00_0018_00_0040_0A54_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a125_1 ( .OUT(na125_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na446_2), .IN5(na2_2), .IN6(1'b0), .IN7(~na436_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x41y34     80'h00_FD00_00_0040_0A31_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a126_1 ( .OUT(na126_1_i), .IN1(1'b1), .IN2(~na7_1), .IN3(1'b1), .IN4(na312_1), .IN5(~na125_1), .IN6(na124_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a126_2 ( .OUT(na126_1), .CLK(~na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na126_1_i) );
// C_ADDF2///ADDF2/      x38y47     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a129_1 ( .OUT(na129_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na151_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a129_4 ( .OUT(na129_2), .COUTY1(na129_4), .IN1(na1_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na151_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y48     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a131_1 ( .OUT(na131_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na93_2),
                     .CINX(1'b0), .CINY1(na129_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a131_4 ( .OUT(na131_2), .COUTY1(na131_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na93_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na93_2), .CINX(1'b0), .CINY1(na129_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y49     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a133_1 ( .OUT(na133_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na36_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na131_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a133_4 ( .OUT(na133_2), .COUTY1(na133_4), .IN1(na36_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na36_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na131_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y50     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a135_1 ( .OUT(na135_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na28_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na133_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a135_4 ( .OUT(na135_2), .COUTY1(na135_4), .IN1(na28_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na28_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na133_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y51     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a137_1 ( .OUT(na137_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na33_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na135_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a137_4 ( .OUT(na137_2), .COUTY1(na137_4), .IN1(na33_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na33_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na135_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y42     80'h00_0078_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na39_2), .IN7(1'b1), .IN8(na59_2),
                     .CINX(1'b0), .CINY1(na152_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a138_4 ( .OUT(na138_2), .COUTY1(na138_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na59_1), .IN5(1'b1), .IN6(na39_2), .IN7(1'b1),
                     .IN8(na59_2), .CINX(1'b0), .CINY1(na152_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y52     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a140_1 ( .OUT(na140_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na29_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na137_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a140_4 ( .OUT(na140_2), .COUTY1(na140_4), .IN1(na29_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na29_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na137_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y53     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a142_1 ( .OUT(na142_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na14_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na140_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a142_4 ( .OUT(na142_2), .IN1(1'b1), .IN2(na14_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na14_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na140_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y43     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a145_1 ( .OUT(na145_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na23_2),
                     .CINX(1'b0), .CINY1(na138_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a145_4 ( .OUT(na145_2), .COUTY1(na145_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na23_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na23_2), .CINX(1'b0), .CINY1(na138_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y44     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a147_1 ( .OUT(na147_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na61_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na145_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a147_4 ( .OUT(na147_2), .COUTY1(na147_4), .IN1(na61_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na61_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na145_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y45     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a149_1 ( .OUT(na149_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na37_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na147_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a149_4 ( .OUT(na149_2), .COUTY1(na149_4), .IN1(na37_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na37_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na147_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y46     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a151_1 ( .OUT(na151_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na41_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na149_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a151_4 ( .OUT(na151_2), .COUTY1(na151_4), .IN1(1'b0), .IN2(1'b0), .IN3(na41_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na41_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na149_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x38y41     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a152_2 ( .OUT(na152_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a152_6 ( .COUTY1(na152_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na152_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x45y37     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a153_1 ( .OUT(na153_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na80_1), .IN7(na79_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na162_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a153_4 ( .OUT(na153_2), .COUTY1(na153_4), .IN1(1'b1), .IN2(na81_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na80_1), .IN7(na79_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na162_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x45y38     80'h00_0078_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a155_1 ( .OUT(na155_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na82_1),
                     .CINX(1'b0), .CINY1(na153_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a155_4 ( .OUT(na155_2), .COUTY1(na155_4), .IN1(1'b0), .IN2(1'b0), .IN3(na83_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na82_1), .CINX(1'b0), .CINY1(na153_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x45y39     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a157_1 ( .OUT(na157_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na84_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na155_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a157_4 ( .OUT(na157_2), .COUTY1(na157_4), .IN1(na85_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na84_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na155_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x45y40     80'h00_0078_00_0020_0C66_0A0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a159_1 ( .OUT(na159_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na86_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na157_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a159_4 ( .OUT(na159_2), .COUTY1(na159_4), .IN1(1'b1), .IN2(na87_1), .IN3(1'b0), .IN4(1'b0), .IN5(na86_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na157_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x45y41     80'h00_0018_00_0010_0666_00A0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a161_1 ( .OUT(na161_1), .IN1(1'b0), .IN2(1'b0), .IN3(na88_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na159_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x45y36     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a162_2 ( .OUT(na162_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a162_6 ( .COUTY1(na162_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na162_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x40y38     80'h00_0078_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a163_1 ( .OUT(na163_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na116_2), .IN7(1'b1), .IN8(na115_2),
                     .CINX(1'b0), .CINY1(na172_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a163_4 ( .OUT(na163_2), .COUTY1(na163_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na115_1), .IN5(1'b1), .IN6(na116_2), .IN7(1'b1),
                     .IN8(na115_2), .CINX(1'b0), .CINY1(na172_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x40y39     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a165_1 ( .OUT(na165_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na103_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na163_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a165_4 ( .OUT(na165_2), .COUTY1(na165_4), .IN1(1'b0), .IN2(1'b0), .IN3(na103_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na103_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na163_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x40y40     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a167_1 ( .OUT(na167_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na90_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na165_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a167_4 ( .OUT(na167_2), .COUTY1(na167_4), .IN1(na90_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na90_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na165_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x40y41     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a169_1 ( .OUT(na169_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na58_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na167_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a169_4 ( .OUT(na169_2), .COUTY1(na169_4), .IN1(1'b0), .IN2(1'b0), .IN3(na58_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na58_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na167_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x40y42     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a171_1 ( .OUT(na171_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na53_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na169_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x40y37     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a172_2 ( .OUT(na172_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a172_6 ( .COUTY1(na172_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na172_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x44y42     80'h00_0078_00_0020_0C66_CC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a173_1 ( .OUT(na173_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na51_1), .IN7(1'b1), .IN8(na443_2),
                     .CINX(1'b0), .CINY1(na182_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a173_4 ( .OUT(na173_2), .COUTY1(na173_4), .IN1(1'b1), .IN2(na47_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na51_1), .IN7(1'b1),
                     .IN8(na443_2), .CINX(1'b0), .CINY1(na182_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x44y43     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a175_1 ( .OUT(na175_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na44_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na173_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a175_4 ( .OUT(na175_2), .COUTY1(na175_4), .IN1(na44_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na44_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na173_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x44y44     80'h00_0078_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a177_1 ( .OUT(na177_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na43_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na175_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a177_4 ( .OUT(na177_2), .COUTY1(na177_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na18_2), .IN5(1'b1), .IN6(na43_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na175_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x44y45     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a179_1 ( .OUT(na179_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na27_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na177_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a179_4 ( .OUT(na179_2), .COUTY1(na179_4), .IN1(na27_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na27_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na177_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x44y46     80'h00_0018_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a181_1 ( .OUT(na181_1), .IN1(1'b1), .IN2(na9_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na179_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x44y41     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a182_2 ( .OUT(na182_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a182_6 ( .COUTY1(na182_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na182_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x44y48     80'h00_0078_00_0020_0C66_CCA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a183_1 ( .OUT(na183_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na447_2), .IN7(1'b1), .IN8(na89_1),
                     .CINX(1'b0), .CINY1(na371_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a183_4 ( .OUT(na183_2), .COUTY1(na183_4), .IN1(1'b0), .IN2(1'b0), .IN3(na52_1), .IN4(1'b1), .IN5(1'b1), .IN6(na447_2), .IN7(1'b1),
                     .IN8(na89_1), .CINX(1'b0), .CINY1(na371_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x44y49     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a185_1 ( .OUT(na185_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na3_2),
                     .CINX(1'b0), .CINY1(na183_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a185_4 ( .OUT(na185_2), .COUTY1(na185_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na3_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na3_2), .CINX(1'b0), .CINY1(na183_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x44y50     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a187_1 ( .OUT(na187_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na101_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na185_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a187_4 ( .OUT(na187_2), .COUTY1(na187_4), .IN1(1'b0), .IN2(1'b0), .IN3(na101_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na101_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na185_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x44y51     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a189_1 ( .OUT(na189_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na100_2),
                     .CINX(1'b0), .CINY1(na187_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a189_4 ( .OUT(na189_2), .COUTY1(na189_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na99_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na100_2), .CINX(1'b0), .CINY1(na187_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x44y52     80'h00_0018_00_0010_0666_00A0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a191_1 ( .OUT(na191_1), .IN1(1'b0), .IN2(1'b0), .IN3(na34_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na189_4), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0014_0016)) 
           _a194 ( .GLB0(na194_1), .GLB1(na194_2), .GLB2(_d0), .GLB3(_d1), .CLK_FB0(_d2), .CLK_FB1(_d3), .CLK_FB2(_d4), .CLK_FB3(_d5),
                   .CLK0_0(na316_6), .CLK0_90(na316_5), .CLK0_180(na316_4), .CLK0_270(na316_3), .CLK0_BYP(1'b0), .CLK1_0(na315_6),
                   .CLK1_90(na315_5), .CLK1_180(na315_4), .CLK1_270(na315_3), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0),
                   .CLK2_270(1'b0), .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0),
                   .USR_GLB0(1'b0), .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0),
                   .USR_FB3(1'b0) );
// C_AND/D///      x34y47     80'h00_FE00_00_0000_0C88_3FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a211_1 ( .OUT(na211_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na21_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a211_2 ( .OUT(na211_1), .CLK(na311_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na211_1_i) );
// C_///AND/D      x35y48     80'h00_FE00_80_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a212_4 ( .OUT(na212_2_i), .IN1(~na67_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a212_5 ( .OUT(na212_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na212_2_i) );
// C_AND/D///      x45y47     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a262_1 ( .OUT(na262_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na34_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a262_2 ( .OUT(na262_1), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na262_1_i) );
// C_///AND/D      x41y44     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a273_4 ( .OUT(na273_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na18_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a273_5 ( .OUT(na273_2), .CLK(na194_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na273_2_i) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a309 ( .Y(na309_1), .I(clk) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a310 ( .Y(na310_1), .I(i_mosi_ILA) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a311 ( .Y(na311_1), .I(i_sclk_ILA) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a312 ( .Y(na312_1), .I(i_ss_ILA) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a313 ( .O(led), .A(na372_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a314 ( .O(o_miso_ILA), .A(na373_10) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_0C_08_0C_20_82)) 
           _a315 ( .USR_PLL_LOCKED_STDY(_d6), .USR_PLL_LOCKED(_d7), .CLK270(na315_3), .CLK180(na315_4), .CLK90(na315_5), .CLK0(na315_6),
                   .CLK_REF_OUT(_d8), .CLK_REF(na322_2), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_3C_08_0C_20_82)) 
           _a316 ( .USR_PLL_LOCKED_STDY(_d9), .USR_PLL_LOCKED(_d10), .CLK270(na316_3), .CLK180(na316_4), .CLK90(na316_5), .CLK0(na316_6),
                   .CLK_REF_OUT(_d11), .CLK_REF(na322_1), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_01_04_05_00_60_00_0D_00_00_00_03_13_00_00_00_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a317 ( .DOA({_d12, _d13, _d14, _d15, _d16, _d17, _d18, _d19, _d20, _d21, _d22, _d23, _d24, _d25, _d26, _d27, _d28, _d29,
                  _d30, _d31, _d32, _d33, _d34, _d35, _d36, _d37, _d38, _d39, _d40, _d41, _d42, _d43, _d44, _d45, _d46, _d47, _d48,
                  _d49, _d50, _d51}),
                   .DOAX({_d52, _d53, _d54, _d55, _d56, _d57, _d58, _d59, _d60, _d61, _d62, _d63, _d64, _d65, _d66, _d67, _d68, _d69,
                  _d70, _d71, _d72, _d73, _d74, _d75, _d76, _d77, _d78, _d79, _d80, _d81, _d82, _d83, _d84, _d85, _d86, _d87, _d88,
                  _d89, _d90, _d91}),
                   .DOB({_d92, _d93, _d94, _d95, _d96, _d97, _d98, _d99, _d100, _d101, _d102, _d103, _d104, _d105, _d106, _d107, _d108,
                  _d109, _d110, _d111, _d112, _d113, _d114, _d115, _d116, _d117, _d118, _d119, _d120, _d121, _d122, _d123, _d124, _d125,
                  _d126, _d127, _d128, _d129, _d130, na317_120}),
                   .DOBX({_d131, _d132, _d133, _d134, _d135, _d136, _d137, _d138, _d139, _d140, _d141, _d142, _d143, _d144, _d145,
                  _d146, _d147, _d148, _d149, _d150, _d151, _d152, _d153, _d154, _d155, _d156, _d157, _d158, _d159, _d160, _d161, _d162,
                  _d163, _d164, _d165, _d166, _d167, _d168, _d169, _d170}),
                   .ECC1B_ERRA({_d171, _d172, _d173, _d174}),
                   .ECC1B_ERRB({_d175, _d176, _d177, _d178}),
                   .ECC2B_ERRA({_d179, _d180, _d181, _d182}),
                   .ECC2B_ERRB({_d183, _d184, _d185, _d186}),
                   .FORW_CAS_WRAO(_d187), .FORW_CAS_WRBO(_d188), .FORW_CAS_BMAO(_d189), .FORW_CAS_BMBO(_d190), .FORW_CAS_RDAO(_d191),
                   .FORW_CAS_RDBO(_d192), .FORW_UADDRAO({_d193, _d194, _d195, _d196, _d197, _d198, _d199, _d200, _d201, _d202, _d203,
                  _d204, _d205, _d206, _d207, _d208}),
                   .FORW_LADDRAO({_d209, _d210, _d211, _d212, _d213, _d214, _d215, _d216, _d217, _d218, _d219, _d220, _d221, _d222,
                  _d223, _d224}),
                   .FORW_UADDRBO({_d225, _d226, _d227, _d228, _d229, _d230, _d231, _d232, _d233, _d234, _d235, _d236, _d237, _d238,
                  _d239, _d240}),
                   .FORW_LADDRBO({_d241, _d242, _d243, _d244, _d245, _d246, _d247, _d248, _d249, _d250, _d251, _d252, _d253, _d254,
                  _d255, _d256}),
                   .FORW_UA0CLKO(_d257), .FORW_UA0ENO(_d258), .FORW_UA0WEO(_d259), .FORW_LA0CLKO(_d260), .FORW_LA0ENO(_d261), .FORW_LA0WEO(_d262),
                   .FORW_UA1CLKO(_d263), .FORW_UA1ENO(_d264), .FORW_UA1WEO(_d265), .FORW_LA1CLKO(_d266), .FORW_LA1ENO(_d267), .FORW_LA1WEO(_d268),
                   .FORW_UB0CLKO(_d269), .FORW_UB0ENO(_d270), .FORW_UB0WEO(_d271), .FORW_LB0CLKO(_d272), .FORW_LB0ENO(_d273), .FORW_LB0WEO(_d274),
                   .FORW_UB1CLKO(_d275), .FORW_UB1ENO(_d276), .FORW_UB1WEO(_d277), .FORW_LB1CLKO(_d278), .FORW_LB1ENO(_d279), .FORW_LB1WEO(_d280),
                   .CLOCKA({_d281, _d282, _d283, _d284}),
                   .CLOCKB({_d285, _d286, _d287, _d288}),
                   .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .CLKB({1'b1, 1'b1, 1'b1, na325_9}),
                   .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .GLWEA({1'b1, 1'b1, 1'b1, na331_10}),
                   .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0({na336_10, na343_9, na346_10, na349_9, na350_10, na360_9, na361_10, na363_9, na365_10, na369_9, na374_10,
                  na375_9, na376_10, na377_9, na378_10, na379_9}),
                   .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB0({na380_10, na381_9, na382_10, na383_9, na384_10, na385_9, na386_10, na387_9, na388_10, na389_9, na390_10,
                  na391_9, na392_10, na393_9, na394_10, na395_9}),
                   .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, na396_10, na397_9, na398_10, na399_9, na400_10, na401_9, na402_10, na403_9, na404_10, na405_9, na406_10,
                  na407_9, na408_10, na409_9, na410_10, na411_9, na412_10, na413_9, na414_10, na415_9}),
                   .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, na416_10, na417_9, na418_10, na419_9, na420_10, na421_9, na422_10, na423_9, na424_10, na425_9, na426_10,
                  na427_9, na428_10, na429_9, na430_10, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .CLOCK1(na194_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                   .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                   .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                   .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                   .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
CC_USR_RSTN            _a318 ( .USR_RSTN(na318_1) );
// C_MX2b////      x43y48     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a319_1 ( .OUT(na319_1), .IN1(1'b1), .IN2(~na25_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na185_2), .IN8(na3_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y37     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a320_1 ( .OUT(na320_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2_1), .IN6(1'b1), .IN7(1'b1), .IN8(na432_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x48y45     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a321_1 ( .OUT(na321_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na446_2), .IN5(1'b0), .IN6(na9_1), .IN7(1'b0), .IN8(na181_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a322 ( .PCLK0(na322_1), .PCLK1(na322_2), .PCLK2(_d289), .PCLK3(_d290), .CLK0(na309_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0),
                   .SER_CLK(1'b0), .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_////RAM_I2      x1y66     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a323_5 ( .OUT(na323_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na318_1), .CP_O(1'b0) );
// C_MX2b////      x41y49     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a324_1 ( .OUT(na324_1), .IN1(1'b1), .IN2(~na25_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na185_1), .IN8(na3_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y33     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a325_1 ( .OUT(na325_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na311_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a325_6 ( .RAM_O1(na325_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na325_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x47y43     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a326_1 ( .OUT(na326_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na446_2), .IN5(na27_1), .IN6(1'b0), .IN7(na179_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x45y42     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a327_1 ( .OUT(na327_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na446_2), .IN5(na27_2), .IN6(1'b0), .IN7(na179_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y43     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a328_1 ( .OUT(na328_1), .IN1(1'b1), .IN2(~na51_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na437_2), .IN8(na177_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x46y41     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a329_1 ( .OUT(na329_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na446_2), .IN5(1'b0), .IN6(na43_1), .IN7(1'b0), .IN8(na177_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x43y40     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a330_1 ( .OUT(na330_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na446_2), .IN5(na44_1), .IN6(1'b0), .IN7(na175_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x27y33     80'h08_0060_00_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a331_4 ( .OUT(na331_2), .IN1(1'b1), .IN2(~na51_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a331_6 ( .RAM_O2(na331_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na331_2), .COMP_OUT(1'b0) );
// C_MX2b////      x42y40     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a332_1 ( .OUT(na332_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na446_2), .IN5(na44_2), .IN6(1'b0), .IN7(na175_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x46y42     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a333_1 ( .OUT(na333_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na446_2), .IN5(1'b0), .IN6(na47_1), .IN7(1'b0), .IN8(na173_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x36y42     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a334_1 ( .OUT(na334_1), .IN1(1'b1), .IN2(na49_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na48_1), .IN8(na68_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x44y40     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a335_1 ( .OUT(na335_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na446_2), .IN5(1'b0), .IN6(na47_2), .IN7(1'b0), .IN8(na173_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a336_4 ( .OUT(na336_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a336_6 ( .RAM_O2(na336_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na336_2), .COMP_OUT(1'b0) );
// C_MX2b////      x43y49     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a337_1 ( .OUT(na337_1), .IN1(1'b1), .IN2(na25_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na52_1), .IN8(na183_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y46     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a338_1 ( .OUT(na338_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na446_2), .IN5(1'b0), .IN6(na9_1), .IN7(1'b0), .IN8(na53_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x33y41     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a339_1 ( .OUT(na339_1), .IN1(na55_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na54_2), .IN6(na63_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y41     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a340_1 ( .OUT(na340_1), .IN1(na55_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na56_1), .IN8(na68_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x40y37     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a341_4 ( .OUT(na341_2), .IN1(1'b0), .IN2(na6_2), .IN3(1'b0), .IN4(na57_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y40     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a342_1 ( .OUT(na342_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na446_2), .IN5(na27_1), .IN6(1'b0), .IN7(na58_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a343_1 ( .OUT(na343_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a343_6 ( .RAM_O1(na343_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na343_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x34y37     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a344_1 ( .OUT(na344_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na446_2), .IN5(na27_2), .IN6(1'b0), .IN7(na58_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x34y35     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a345_1 ( .OUT(na345_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na446_2), .IN5(1'b0), .IN6(na51_1), .IN7(1'b0), .IN8(na115_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y39     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a346_4 ( .OUT(na346_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na53_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a346_6 ( .RAM_O2(na346_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na346_2), .COMP_OUT(1'b0) );
// C_MX2b////      x42y46     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a347_1 ( .OUT(na347_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na446_2), .IN5(1'b0), .IN6(na451_2), .IN7(1'b0), .IN8(na18_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x36y37     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a348_1 ( .OUT(na348_1), .IN1(1'b1), .IN2(~na51_2), .IN3(1'b0), .IN4(1'b0), .IN5(na90_2), .IN6(na43_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y39     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a349_1 ( .OUT(na349_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na58_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a349_6 ( .RAM_O1(na349_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na349_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y38     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a350_4 ( .OUT(na350_2), .IN1(1'b1), .IN2(1'b1), .IN3(na58_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a350_6 ( .RAM_O2(na350_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na350_2), .COMP_OUT(1'b0) );
// C_MX2b////      x34y42     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a351_1 ( .OUT(na351_1), .IN1(~na55_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na40_1), .IN6(na97_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y49     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a352_1 ( .OUT(na352_1), .IN1(1'b1), .IN2(na25_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na34_2), .IN8(na191_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x45y49     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a353_1 ( .OUT(na353_1), .IN1(1'b1), .IN2(~na25_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na189_2), .IN8(na99_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x46y47     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a354_1 ( .OUT(na354_1), .IN1(1'b1), .IN2(~na25_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na189_1), .IN8(na100_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x41y48     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a355_1 ( .OUT(na355_1), .IN1(1'b1), .IN2(na25_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na101_1), .IN8(na187_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y50     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a356_1 ( .OUT(na356_1), .IN1(1'b1), .IN2(na25_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na101_2), .IN8(na187_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y42     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a357_1 ( .OUT(na357_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na446_2), .IN5(na44_1), .IN6(1'b0), .IN7(na103_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x34y43     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a358_1 ( .OUT(na358_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na446_2), .IN5(na44_2), .IN6(1'b0), .IN7(na103_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x36y47     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a359_1 ( .OUT(na359_1), .IN1(1'b1), .IN2(~na49_2), .IN3(1'b0), .IN4(1'b0), .IN5(na40_1), .IN6(na105_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y38     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a360_1 ( .OUT(na360_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na90_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a360_6 ( .RAM_O1(na360_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na360_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y37     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a361_4 ( .OUT(na361_2), .IN1(na90_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a361_6 ( .RAM_O2(na361_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na361_2), .COMP_OUT(1'b0) );
// C_MX2b////      x45y46     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a362_1 ( .OUT(na362_1), .IN1(1'b1), .IN2(na25_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na52_2), .IN8(na183_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y37     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a363_1 ( .OUT(na363_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na103_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a363_6 ( .RAM_O1(na363_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na363_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x39y40     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a364_1 ( .OUT(na364_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na6_2), .IN7(na107_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y36     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a365_4 ( .OUT(na365_2), .IN1(1'b1), .IN2(1'b1), .IN3(na103_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a365_6 ( .RAM_O2(na365_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na365_2), .COMP_OUT(1'b0) );
// C_MX2b////      x34y46     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a366_1 ( .OUT(na366_1), .IN1(~na114_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na16_2), .IN6(na13_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x44y37     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a367_1 ( .OUT(na367_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na446_2), .IN5(1'b0), .IN6(na47_1), .IN7(1'b0), .IN8(na115_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x33y42     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a368_1 ( .OUT(na368_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na446_2), .IN5(1'b0), .IN6(na116_2), .IN7(1'b0), .IN8(na443_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a369_1 ( .OUT(na369_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a369_6 ( .RAM_O1(na369_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na369_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x34y45     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a370_1 ( .OUT(na370_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2_2), .IN6(1'b1), .IN7(na107_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x44y47     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a371_2 ( .OUT(na371_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a371_6 ( .COUTY1(na371_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na371_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x107y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a372_4 ( .OUT(na372_2), .IN1(1'b1), .IN2(na14_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a372_6 ( .RAM_O2(na372_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na372_2), .COMP_OUT(1'b0) );
// C_///AND/      x19y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a373_4 ( .OUT(na373_2), .IN1(1'b1), .IN2(na126_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a373_6 ( .RAM_O2(na373_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na373_2), .COMP_OUT(1'b0) );
// C_///AND/      x28y35     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a374_4 ( .OUT(na374_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na115_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a374_6 ( .RAM_O2(na374_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na374_2), .COMP_OUT(1'b0) );
// C_AND////      x28y35     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a375_1 ( .OUT(na375_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na116_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a375_6 ( .RAM_O1(na375_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na375_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y34     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a376_4 ( .OUT(na376_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na115_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a376_6 ( .RAM_O2(na376_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na376_2), .COMP_OUT(1'b0) );
// C_AND////      x28y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a377_1 ( .OUT(na377_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a377_6 ( .RAM_O1(na377_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na377_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a378_4 ( .OUT(na378_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a378_6 ( .RAM_O2(na378_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na378_2), .COMP_OUT(1'b0) );
// C_AND////      x28y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a379_1 ( .OUT(na379_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a379_6 ( .RAM_O1(na379_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na379_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a380_4 ( .OUT(na380_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a380_6 ( .RAM_O2(na380_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na380_2), .COMP_OUT(1'b0) );
// C_AND////      x37y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a381_1 ( .OUT(na381_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a381_6 ( .RAM_O1(na381_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na381_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y39     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a382_4 ( .OUT(na382_2), .IN1(1'b1), .IN2(1'b1), .IN3(na88_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a382_6 ( .RAM_O2(na382_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na382_2), .COMP_OUT(1'b0) );
// C_AND////      x37y39     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a383_1 ( .OUT(na383_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na87_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a383_6 ( .RAM_O1(na383_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na383_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y38     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a384_4 ( .OUT(na384_2), .IN1(na86_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a384_6 ( .RAM_O2(na384_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na384_2), .COMP_OUT(1'b0) );
// C_AND////      x37y38     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a385_1 ( .OUT(na385_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na85_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a385_6 ( .RAM_O1(na385_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na385_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y37     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a386_4 ( .OUT(na386_2), .IN1(na84_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a386_6 ( .RAM_O2(na386_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na386_2), .COMP_OUT(1'b0) );
// C_AND////      x37y37     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a387_1 ( .OUT(na387_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na83_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a387_6 ( .RAM_O1(na387_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na387_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y36     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a388_4 ( .OUT(na388_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na82_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a388_6 ( .RAM_O2(na388_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na388_2), .COMP_OUT(1'b0) );
// C_AND////      x37y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a389_1 ( .OUT(na389_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a389_6 ( .RAM_O1(na389_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na389_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y35     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a390_4 ( .OUT(na390_2), .IN1(1'b1), .IN2(na81_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a390_6 ( .RAM_O2(na390_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na390_2), .COMP_OUT(1'b0) );
// C_AND////      x37y35     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a391_1 ( .OUT(na391_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na80_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a391_6 ( .RAM_O1(na391_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na391_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y34     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a392_4 ( .OUT(na392_2), .IN1(1'b1), .IN2(1'b1), .IN3(na79_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a392_6 ( .RAM_O2(na392_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na392_2), .COMP_OUT(1'b0) );
// C_AND////      x37y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a393_1 ( .OUT(na393_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a393_6 ( .RAM_O1(na393_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na393_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a394_4 ( .OUT(na394_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a394_6 ( .RAM_O2(na394_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na394_2), .COMP_OUT(1'b0) );
// C_AND////      x37y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a395_1 ( .OUT(na395_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a395_6 ( .RAM_O1(na395_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na395_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a396_4 ( .OUT(na396_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a396_6 ( .RAM_O2(na396_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na396_2), .COMP_OUT(1'b0) );
// C_AND////      x30y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a397_1 ( .OUT(na397_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a397_6 ( .RAM_O1(na397_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na397_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a398_4 ( .OUT(na398_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a398_6 ( .RAM_O2(na398_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na398_2), .COMP_OUT(1'b0) );
// C_AND////      x30y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a399_1 ( .OUT(na399_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a399_6 ( .RAM_O1(na399_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na399_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a400_4 ( .OUT(na400_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a400_6 ( .RAM_O2(na400_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na400_2), .COMP_OUT(1'b0) );
// C_AND////      x32y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a401_1 ( .OUT(na401_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a401_6 ( .RAM_O1(na401_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na401_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a402_4 ( .OUT(na402_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a402_6 ( .RAM_O2(na402_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na402_2), .COMP_OUT(1'b0) );
// C_AND////      x32y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a403_1 ( .OUT(na403_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a403_6 ( .RAM_O1(na403_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na403_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y38     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a404_4 ( .OUT(na404_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a404_6 ( .RAM_O2(na404_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na404_2), .COMP_OUT(1'b0) );
// C_AND////      x32y38     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a405_1 ( .OUT(na405_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a405_6 ( .RAM_O1(na405_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na405_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y37     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a406_4 ( .OUT(na406_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a406_6 ( .RAM_O2(na406_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na406_2), .COMP_OUT(1'b0) );
// C_AND////      x32y37     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a407_1 ( .OUT(na407_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a407_6 ( .RAM_O1(na407_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na407_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y36     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a408_4 ( .OUT(na408_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a408_6 ( .RAM_O2(na408_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na408_2), .COMP_OUT(1'b0) );
// C_AND////      x32y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a409_1 ( .OUT(na409_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a409_6 ( .RAM_O1(na409_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na409_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y35     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a410_4 ( .OUT(na410_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a410_6 ( .RAM_O2(na410_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na410_2), .COMP_OUT(1'b0) );
// C_AND////      x32y35     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a411_1 ( .OUT(na411_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a411_6 ( .RAM_O1(na411_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na411_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y34     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a412_4 ( .OUT(na412_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a412_6 ( .RAM_O2(na412_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na412_2), .COMP_OUT(1'b0) );
// C_AND////      x32y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a413_1 ( .OUT(na413_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a413_6 ( .RAM_O1(na413_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na413_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a414_4 ( .OUT(na414_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a414_6 ( .RAM_O2(na414_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na414_2), .COMP_OUT(1'b0) );
// C_AND////      x32y33     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a415_1 ( .OUT(na415_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na309_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a415_6 ( .RAM_O1(na415_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na415_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a416_4 ( .OUT(na416_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a416_6 ( .RAM_O2(na416_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na416_2), .COMP_OUT(1'b0) );
// C_AND////      x29y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a417_1 ( .OUT(na417_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a417_6 ( .RAM_O1(na417_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na417_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a418_4 ( .OUT(na418_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a418_6 ( .RAM_O2(na418_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na418_2), .COMP_OUT(1'b0) );
// C_AND////      x29y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a419_1 ( .OUT(na419_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a419_6 ( .RAM_O1(na419_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na419_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a420_4 ( .OUT(na420_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a420_6 ( .RAM_O2(na420_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na420_2), .COMP_OUT(1'b0) );
// C_AND////      x31y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a421_1 ( .OUT(na421_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a421_6 ( .RAM_O1(na421_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na421_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a422_4 ( .OUT(na422_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a422_6 ( .RAM_O2(na422_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na422_2), .COMP_OUT(1'b0) );
// C_AND////      x31y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a423_1 ( .OUT(na423_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a423_6 ( .RAM_O1(na423_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na423_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y38     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a424_4 ( .OUT(na424_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a424_6 ( .RAM_O2(na424_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na424_2), .COMP_OUT(1'b0) );
// C_AND////      x31y38     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a425_1 ( .OUT(na425_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a425_6 ( .RAM_O1(na425_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na425_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y37     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a426_4 ( .OUT(na426_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a426_6 ( .RAM_O2(na426_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na426_2), .COMP_OUT(1'b0) );
// C_AND////      x31y37     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a427_1 ( .OUT(na427_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a427_6 ( .RAM_O1(na427_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na427_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y36     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a428_4 ( .OUT(na428_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a428_6 ( .RAM_O2(na428_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na428_2), .COMP_OUT(1'b0) );
// C_AND////      x31y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a429_1 ( .OUT(na429_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a429_6 ( .RAM_O1(na429_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na429_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y35     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a430_4 ( .OUT(na430_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a430_6 ( .RAM_O2(na430_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na430_2), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x34y33     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a431_2 ( .OUT(na431_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na317_120), .CP_O(1'b0) );
// C_////Bridge      x36y36     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a432_5 ( .OUT(na432_2), .IN1(na2_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y38     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a433_5 ( .OUT(na433_2), .IN1(1'b0), .IN2(na6_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y35     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a434_5 ( .OUT(na434_2), .IN1(1'b0), .IN2(na10_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y48     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a435_5 ( .OUT(na435_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na16_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y35     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a436_5 ( .OUT(na436_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na17_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y41     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a437_5 ( .OUT(na437_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na18_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y43     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a438_5 ( .OUT(na438_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na21_1) );
// C_////Bridge      x46y45     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a439_5 ( .OUT(na439_2), .IN1(1'b0), .IN2(na25_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y46     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a440_5 ( .OUT(na440_2), .IN1(1'b0), .IN2(na25_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y47     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a441_5 ( .OUT(na441_2), .IN1(1'b0), .IN2(na25_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y38     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a442_5 ( .OUT(na442_2), .IN1(1'b0), .IN2(1'b0), .IN3(na45_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y40     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a443_5 ( .OUT(na443_2), .IN1(1'b0), .IN2(na47_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y42     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a444_5 ( .OUT(na444_2), .IN1(1'b0), .IN2(na51_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y43     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a445_5 ( .OUT(na445_2), .IN1(1'b0), .IN2(na51_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y42     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a446_5 ( .OUT(na446_2), .IN1(1'b0), .IN2(na51_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y48     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a447_5 ( .OUT(na447_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na52_2), .IN8(1'b0) );
// C_////Bridge      x41y35     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a448_5 ( .OUT(na448_2), .IN1(1'b0), .IN2(na66_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y33     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a449_5 ( .OUT(na449_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na66_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y49     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a450_5 ( .OUT(na450_2), .IN1(na67_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y44     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a451_5 ( .OUT(na451_2), .IN1(na90_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y46     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a452_5 ( .OUT(na452_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na106_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y34     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a453_5 ( .OUT(na453_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na163_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y36     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a454_5 ( .OUT(na454_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na163_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y35     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a455_5 ( .OUT(na455_2), .IN1(1'b0), .IN2(1'b0), .IN3(na165_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y37     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a456_5 ( .OUT(na456_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na165_2), .IN8(1'b0) );
// C_////Bridge      x41y38     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a457_5 ( .OUT(na457_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na167_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y36     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a458_5 ( .OUT(na458_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na167_2) );
// C_////Bridge      x43y39     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a459_5 ( .OUT(na459_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na169_1), .IN8(1'b0) );
// C_////Bridge      x41y37     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a460_5 ( .OUT(na460_2), .IN1(1'b0), .IN2(1'b0), .IN3(na169_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y38     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a461_5 ( .OUT(na461_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na171_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
endmodule
