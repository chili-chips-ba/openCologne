//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 September 2024)
//  Compile Time: 2024-09-03 10:56:35
//  Program Run:  2024-09-23 19:15:20
//  Program Call: /home/user/FPGA/Boards/GateMate/cc-toolchain-linux//bin/p_r/p_r -v -i net/top_synth.v -o top -ccf top.ccf -cCP 
//  File Type:    Verilog

// Gatecount:    683
module top (arst_n , clk , uart_rx_serial ,
       bck , clk_check , din , led , lrck 
       ) ;

input  arst_n;
input  clk;
input  uart_rx_serial;

output bck;
output clk_check;
output din;
output [7:0]led;
output lrck;



wire [7:0]led;
wire bck;
wire clk;
wire din;
wire lrck;
wire na1_1;
wire na1_1_i;
wire na3_1;
wire na3_2;
wire na4_2;
wire na7_1;
wire na7_2;
wire na8_1;
wire na8_2;
wire na9_2;
wire arst_n;
wire na10_1;
wire na10_2;
wire na12_1;
wire na12_1_i;
wire na13_1;
wire na13_2;
wire na15_1;
wire na17_1;
wire na18_1;
wire na22_1;
wire na22_2;
wire na23_1;
wire na23_1_i;
wire na27_1;
wire na27_1_i;
wire na30_1;
wire na30_1_i;
wire na33_1;
wire na33_1_i;
wire na36_1;
wire na36_1_i;
wire na37_2;
wire na41_1;
wire na41_1_i;
wire na42_2;
wire na43_1;
wire na43_2;
wire na46_1;
wire na46_1_i;
wire na48_1;
wire na49_2;
wire na50_1;
wire na50_1_i;
wire na53_1;
wire na54_1;
wire na54_1_i;
wire na56_1;
wire na57_1;
wire na59_1;
wire na59_1_i;
wire na62_1;
wire na62_1_i;
wire na64_2;
wire na65_1;
wire na66_1;
wire na66_1_i;
wire na69_1;
wire na69_1_i;
wire na72_1;
wire na72_1_i;
wire na75_1;
wire na75_1_i;
wire na78_1;
wire na78_1_i;
wire na81_1;
wire na81_1_i;
wire na84_1;
wire na84_1_i;
wire na87_1;
wire na87_1_i;
wire na90_1;
wire na90_1_i;
wire na93_1;
wire na93_1_i;
wire na96_1;
wire na96_1_i;
wire na99_1;
wire na99_1_i;
wire na102_1;
wire na102_1_i;
wire na105_1;
wire na105_1_i;
wire na107_2;
wire na109_1;
wire na109_1_i;
wire na112_1;
wire na112_1_i;
wire na115_1;
wire na115_1_i;
wire na117_1;
wire na119_1;
wire na119_1_i;
wire na122_1;
wire na122_1_i;
wire na125_1;
wire na125_1_i;
wire na128_1;
wire na128_1_i;
wire na131_1;
wire na131_1_i;
wire na134_1;
wire na134_1_i;
wire na137_1;
wire na137_1_i;
wire na138_1;
wire na138_2;
wire na141_1;
wire na141_1_i;
wire na145_2;
wire na146_1;
wire na146_1_i;
wire na149_1;
wire na149_1_i;
wire na152_1;
wire na152_1_i;
wire na155_1;
wire na155_1_i;
wire na158_1;
wire na158_1_i;
wire na161_1;
wire na161_1_i;
wire na164_1;
wire na164_1_i;
wire na167_1;
wire na167_1_i;
wire na170_1;
wire na170_1_i;
wire na173_1;
wire na173_1_i;
wire na176_1;
wire na176_1_i;
wire na179_1;
wire na179_1_i;
wire na182_1;
wire na182_1_i;
wire na186_1;
wire na186_1_i;
wire na189_1;
wire na189_1_i;
wire na191_1;
wire na192_2;
wire na193_1;
wire na193_1_i;
wire na196_1;
wire na196_1_i;
wire na199_1;
wire na199_1_i;
wire na202_1;
wire na202_1_i;
wire na205_1;
wire na205_1_i;
wire na209_1;
wire na209_1_i;
wire na212_1;
wire na212_1_i;
wire na215_1;
wire na215_1_i;
wire na218_1;
wire na218_1_i;
wire na221_1;
wire na221_1_i;
wire na224_1;
wire na224_1_i;
wire na227_1;
wire na229_1;
wire na230_2;
wire na231_1;
wire na232_1;
wire na233_1;
wire na233_2;
wire na234_1;
wire na235_2;
wire na236_1;
wire na236_1_i;
wire na237_1;
wire na237_1_i;
wire na237_2;
wire na237_2_i;
wire na239_1;
wire na239_1_i;
wire na239_2;
wire na239_2_i;
wire na241_1;
wire na241_1_i;
wire na241_2;
wire na241_2_i;
wire na243_1;
wire na243_1_i;
wire na243_2;
wire na243_2_i;
wire na245_1;
wire na245_1_i;
wire na245_2;
wire na245_2_i;
wire na246_2;
wire na246_2_i;
wire na247_1;
wire na247_1_i;
wire na247_2;
wire na247_2_i;
wire na249_2;
wire na249_2_i;
wire na250_2;
wire na250_2_i;
wire na251_1;
wire na251_1_i;
wire na252_1;
wire na253_2;
wire na254_1;
wire na257_1;
wire na257_2;
wire na258_1;
wire na258_1_i;
wire na259_1;
wire na260_1;
wire na260_2;
wire na261_2;
wire na262_1;
wire na262_1_i;
wire na263_1;
wire na265_1;
wire na265_1_i;
wire na265_2;
wire na265_2_i;
wire na266_2;
wire na267_1;
wire na268_1;
wire na269_1;
wire na270_2;
wire na271_1;
wire na271_1_i;
wire na271_2;
wire na271_2_i;
wire na272_1;
wire na272_1_i;
wire na273_1;
wire na274_1;
wire na274_1_i;
wire na275_2;
wire na276_1;
wire na276_1_i;
wire na277_1;
wire na278_1;
wire na278_1_i;
wire na279_2;
wire na280_1;
wire na280_1_i;
wire na281_2;
wire na282_1;
wire na282_1_i;
wire na283_1;
wire na283_1_i;
wire na284_1;
wire na284_1_i;
wire na315_1;
wire na315_1_i;
wire na318_4;
wire na320_4;
wire na322_4;
wire na323_4;
wire na325_4;
wire na327_4;
wire na329_4;
wire na331_4;
wire na332_1;
wire na332_4;
wire na334_1;
wire na334_2;
wire na334_4;
wire na336_1;
wire na336_2;
wire na336_4;
wire na338_1;
wire na338_2;
wire na338_4;
wire na340_1;
wire na340_2;
wire na340_4;
wire na342_1;
wire na342_2;
wire na342_4;
wire na343_1;
wire na343_2;
wire na343_4;
wire na345_1;
wire na345_2;
wire na345_4;
wire na347_1;
wire na347_2;
wire na347_4;
wire na349_1;
wire na349_2;
wire na349_4;
wire na351_1;
wire na351_2;
wire na351_4;
wire na353_1;
wire na353_2;
wire na353_4;
wire na356_1;
wire na356_2;
wire na356_4;
wire na358_1;
wire na358_2;
wire na358_4;
wire na360_1;
wire na360_2;
wire na360_4;
wire na362_1;
wire na362_2;
wire na362_4;
wire na364_1;
wire na364_2;
wire na364_4;
wire na365_1;
wire na365_2;
wire na365_4;
wire na367_1;
wire na367_2;
wire na367_4;
wire na369_1;
wire na369_2;
wire na369_4;
wire na371_1;
wire na371_2;
wire na371_4;
wire na373_1;
wire na373_2;
wire na373_4;
wire na375_1;
wire na375_2;
wire na375_4;
wire na378_1;
wire na378_2;
wire na378_4;
wire na380_1;
wire na380_2;
wire na380_4;
wire na382_1;
wire na382_2;
wire na382_4;
wire na384_1;
wire na384_2;
wire na384_4;
wire na386_1;
wire na386_2;
wire na386_4;
wire na387_1;
wire na387_2;
wire na387_4;
wire na389_1;
wire na389_2;
wire na392_1;
wire na392_2;
wire na392_4;
wire na394_1;
wire na394_2;
wire na394_4;
wire na395_1;
wire na395_4;
wire na397_1;
wire na397_2;
wire na397_4;
wire na399_1;
wire na399_2;
wire na399_4;
wire na401_1;
wire na401_2;
wire na401_4;
wire na403_1;
wire na403_2;
wire na403_4;
wire na405_1;
wire na405_2;
wire na405_4;
wire na406_1;
wire na406_2;
wire na406_4;
wire na408_1;
wire na408_2;
wire na408_4;
wire na410_1;
wire na410_2;
wire na410_4;
wire na412_1;
wire na412_2;
wire na412_4;
wire na414_1;
wire na414_2;
wire na414_4;
wire na416_1;
wire na416_2;
wire na416_4;
wire na419_1;
wire na419_2;
wire na419_4;
wire na421_1;
wire na421_2;
wire na421_4;
wire na423_1;
wire na423_2;
wire na423_4;
wire na425_1;
wire na425_2;
wire na425_4;
wire na427_1;
wire na427_2;
wire na427_4;
wire na428_1;
wire na428_2;
wire na428_4;
wire na430_1;
wire na430_2;
wire na430_4;
wire na432_1;
wire na432_2;
wire na432_4;
wire na434_1;
wire na434_2;
wire na434_4;
wire na436_1;
wire na436_2;
wire na436_4;
wire na438_1;
wire na438_2;
wire na438_4;
wire na441_1;
wire na441_2;
wire na441_4;
wire na443_1;
wire na443_2;
wire na443_4;
wire na445_1;
wire na445_2;
wire na445_4;
wire na447_1;
wire na447_2;
wire na447_4;
wire na449_1;
wire na449_2;
wire na449_4;
wire na450_1;
wire na450_2;
wire na450_4;
wire na452_1;
wire na452_2;
wire na452_4;
wire na454_1;
wire na456_1;
wire na456_2;
wire na456_4;
wire na458_1;
wire na458_2;
wire na458_4;
wire na459_1;
wire na459_4;
wire na460_1;
wire na460_1_i;
wire na460_2;
wire na462_1;
wire na462_4;
wire na463_1;
wire na463_1_i;
wire na463_2;
wire na463_4;
wire na465_1;
wire na465_1_i;
wire na465_2;
wire na465_4;
wire na467_1;
wire na467_1_i;
wire na468_1;
wire na468_1_i;
wire na468_2;
wire na468_4;
wire na469_1;
wire na469_1_i;
wire na469_2;
wire na469_4;
wire na471_1;
wire na471_1_i;
wire na471_2;
wire na471_4;
wire na473_1;
wire na473_1_i;
wire na473_2;
wire na473_4;
wire na475_1;
wire na475_1_i;
wire na475_2;
wire na475_4;
wire na477_1;
wire na477_1_i;
wire na477_2;
wire na477_4;
wire na480_1;
wire na480_1_i;
wire na480_2;
wire na480_4;
wire na482_1;
wire na482_1_i;
wire na482_2;
wire na482_4;
wire na484_1;
wire na484_1_i;
wire na484_2;
wire na484_4;
wire na486_1;
wire na486_1_i;
wire na486_2;
wire na486_4;
wire na488_1;
wire na488_1_i;
wire na488_2;
wire na488_4;
wire na490_1;
wire na490_1_i;
wire na490_2;
wire na490_4;
wire na491_1;
wire na491_1_i;
wire na491_2;
wire na491_4;
wire na493_1;
wire na493_1_i;
wire na493_2;
wire na493_4;
wire na495_1;
wire na495_1_i;
wire na495_2;
wire na495_4;
wire na497_1;
wire na497_1_i;
wire na497_2;
wire na497_4;
wire na499_1;
wire na499_1_i;
wire na499_2;
wire na499_4;
wire na502_1;
wire na502_1_i;
wire na502_2;
wire na502_4;
wire na504_1;
wire na504_1_i;
wire na504_2;
wire na504_4;
wire na506_1;
wire na506_1_i;
wire na506_2;
wire na506_4;
wire na508_1;
wire na508_1_i;
wire na508_2;
wire na508_4;
wire na510_1;
wire na510_1_i;
wire na510_2;
wire na510_4;
wire na512_1;
wire na512_1_i;
wire na512_2;
wire na512_4;
wire na513_1;
wire na513_1_i;
wire na513_2;
wire na513_4;
wire na515_1;
wire na515_1_i;
wire na515_2;
wire na515_4;
wire na517_1;
wire na517_1_i;
wire na517_2;
wire na517_4;
wire na519_1;
wire na519_1_i;
wire na519_2;
wire na519_4;
wire na521_1;
wire na521_1_i;
wire na521_2;
wire na521_4;
wire na524_1;
wire na524_1_i;
wire na524_2;
wire na524_4;
wire na526_1;
wire na526_1_i;
wire na526_2;
wire na528_1;
wire na528_1_i;
wire na528_2;
wire na528_4;
wire na530_1;
wire na530_1_i;
wire na530_2;
wire na530_4;
wire na532_1;
wire na532_4;
wire na533_1;
wire na533_2;
wire na535_1;
wire na535_4;
wire na537_1;
wire na537_2;
wire na537_4;
wire na539_1;
wire na539_2;
wire na539_4;
wire na541_1;
wire na542_1;
wire na542_2;
wire na542_4;
wire na544_1;
wire na544_2;
wire na544_4;
wire na546_1;
wire na546_2;
wire na546_4;
wire na548_1;
wire na548_2;
wire na548_4;
wire na550_1;
wire na550_2;
wire na550_4;
wire na551_1;
wire na551_4;
wire na552_1;
wire na552_2;
wire na552_4;
wire na554_1;
wire na554_4;
wire na555_1;
wire na555_4;
wire na557_1;
wire na557_2;
wire na557_4;
wire na559_1;
wire na559_2;
wire na559_4;
wire na561_1;
wire na561_2;
wire na561_4;
wire na563_1;
wire na563_2;
wire na563_4;
wire na565_1;
wire na565_2;
wire na565_4;
wire na566_1;
wire na566_2;
wire na566_4;
wire na568_1;
wire na568_2;
wire na568_4;
wire na570_1;
wire na570_2;
wire na570_4;
wire na572_1;
wire na572_2;
wire na572_4;
wire na574_1;
wire na574_2;
wire na574_4;
wire na576_1;
wire na576_2;
wire na576_4;
wire na579_1;
wire na579_2;
wire na579_4;
wire na581_1;
wire na581_2;
wire na581_4;
wire na583_1;
wire na583_2;
wire na583_4;
wire na585_1;
wire na585_2;
wire na585_4;
wire na587_1;
wire na587_2;
wire na587_4;
wire na588_1;
wire na588_2;
wire na588_4;
wire na590_1;
wire na590_2;
wire na590_4;
wire na592_1;
wire na592_2;
wire na592_4;
wire na594_1;
wire na594_2;
wire na594_4;
wire na596_1;
wire na596_2;
wire na596_4;
wire na598_1;
wire na598_2;
wire na598_4;
wire na601_1;
wire na601_2;
wire na601_4;
wire na603_1;
wire na603_2;
wire na603_4;
wire na605_1;
wire na605_2;
wire na605_4;
wire na607_1;
wire na607_2;
wire na607_4;
wire na609_1;
wire na609_2;
wire na609_4;
wire na610_1;
wire na610_2;
wire na610_4;
wire na612_1;
wire na612_2;
wire na615_1;
wire na615_2;
wire na615_4;
wire na617_1;
wire na617_2;
wire na617_4;
wire na618_1;
wire na618_4;
wire na620_1;
wire na620_2;
wire na620_4;
wire na622_1;
wire na622_2;
wire na622_4;
wire na624_1;
wire na624_2;
wire na624_4;
wire na626_1;
wire na626_2;
wire na626_4;
wire na628_1;
wire na628_2;
wire na628_4;
wire na629_1;
wire na629_2;
wire na629_4;
wire na631_1;
wire na631_2;
wire na631_4;
wire na633_1;
wire na633_2;
wire na633_4;
wire na635_1;
wire na635_2;
wire na635_4;
wire na637_1;
wire na637_2;
wire na637_4;
wire na639_1;
wire na639_2;
wire na639_4;
wire na642_1;
wire na642_2;
wire na642_4;
wire na644_1;
wire na644_2;
wire na644_4;
wire na646_1;
wire na646_2;
wire na646_4;
wire na648_1;
wire na648_2;
wire na648_4;
wire na650_1;
wire na650_2;
wire na650_4;
wire na651_1;
wire na651_2;
wire na651_4;
wire na653_1;
wire na653_2;
wire na653_4;
wire na655_1;
wire na655_2;
wire na655_4;
wire na657_1;
wire na657_2;
wire na657_4;
wire na659_1;
wire na659_2;
wire na659_4;
wire na661_1;
wire na661_2;
wire na661_4;
wire na664_1;
wire na664_2;
wire na664_4;
wire na666_1;
wire na666_2;
wire na666_4;
wire na668_1;
wire na668_2;
wire na668_4;
wire na670_1;
wire na670_2;
wire na670_4;
wire na672_1;
wire na672_2;
wire na672_4;
wire na673_1;
wire na673_2;
wire na673_4;
wire na675_1;
wire na675_2;
wire na675_4;
wire na677_1;
wire na679_1;
wire na679_2;
wire na679_4;
wire na681_1;
wire na681_2;
wire na681_4;
wire na685_1;
wire na685_2;
wire na685_3;
wire na703_1;
wire na703_1_i;
wire na703_2;
wire na703_2_i;
wire na704_1;
wire na704_1_i;
wire na704_2;
wire na704_2_i;
wire na707_2;
wire na707_2_i;
wire na708_1;
wire na708_1_i;
wire na709_1;
wire na709_1_i;
wire na710_1;
wire na710_1_i;
wire na717_2;
wire na717_2_i;
wire na719_1;
wire na719_1_i;
wire na721_2;
wire na721_2_i;
wire na723_2;
wire na723_2_i;
wire na725_2;
wire na725_2_i;
wire na727_1;
wire na727_1_i;
wire na729_2;
wire na729_2_i;
wire na731_1;
wire na731_1_i;
wire na733_1;
wire na733_1_i;
wire na735_1;
wire na735_1_i;
wire na737_2;
wire na737_2_i;
wire na739_1;
wire na739_1_i;
wire na741_2;
wire na741_2_i;
wire na743_2;
wire na743_2_i;
wire na745_2;
wire na745_2_i;
wire na747_1;
wire na747_1_i;
wire na749_1;
wire na749_1_i;
wire na751_1;
wire na751_1_i;
wire na753_2;
wire na753_2_i;
wire na755_2;
wire na755_2_i;
wire na757_2;
wire na757_2_i;
wire na759_1;
wire na759_1_i;
wire na761_2;
wire na761_2_i;
wire na763_1;
wire na763_1_i;
wire na765_1;
wire na765_1_i;
wire na767_1;
wire na767_1_i;
wire na769_2;
wire na769_2_i;
wire na771_1;
wire na771_1_i;
wire na773_2;
wire na773_2_i;
wire na775_2;
wire na775_2_i;
wire na777_2;
wire na777_2_i;
wire na779_1;
wire na779_1_i;
wire na780_1;
wire na780_1_i;
wire na780_2;
wire na780_2_i;
wire na782_2;
wire na782_2_i;
wire na784_1;
wire na784_1_i;
wire na788_1;
wire na788_1_i;
wire na789_1;
wire na789_1_i;
wire na791_2;
wire na791_2_i;
wire na857_1;
wire na857_1_i;
wire na857_2;
wire na857_2_i;
wire na869_1;
wire na870_1;
wire na871_1;
wire na872_1;
wire na873_1;
wire na874_1;
wire na875_1;
wire na876_1;
wire na877_1;
wire na878_1;
wire na880_1;
wire na882_1;
wire na894_1;
wire na895_3;
wire na895_4;
wire na895_5;
wire na895_6;
wire na896_2;
wire na896_2_i;
wire na897_1;
wire na897_9;
wire na898_1;
wire na898_4;
wire na899_1;
wire na900_1;
wire na901_1;
wire na902_1;
wire na902_2;
wire na903_2;
wire na904_1;
wire na904_9;
wire na905_2;
wire na906_1;
wire na907_1;
wire na907_9;
wire na908_2;
wire na909_1;
wire na909_9;
wire na910_2;
wire na911_1;
wire na911_9;
wire na912_1;
wire na913_1;
wire na913_2;
wire na914_2;
wire na915_2;
wire na916_1;
wire na917_1;
wire na917_9;
wire na918_2;
wire na919_1;
wire na920_1;
wire na920_2;
wire na921_1;
wire na922_1;
wire na922_9;
wire na923_2;
wire na924_2;
wire na925_1;
wire na925_2;
wire na926_2;
wire na927_1;
wire na927_2;
wire na928_1;
wire na928_9;
wire na929_2;
wire na930_1;
wire na930_2;
wire na931_1;
wire na932_1;
wire na932_9;
wire na933_2;
wire na934_2;
wire na935_1;
wire na935_9;
wire na936_1;
wire na937_2;
wire na938_1;
wire na938_2;
wire na939_2;
wire na940_1;
wire na940_9;
wire na941_1;
wire na941_2;
wire na942_1;
wire na943_1;
wire na943_9;
wire na944_2;
wire na945_1;
wire na945_2;
wire na946_1;
wire na946_9;
wire na947_2;
wire na948_1;
wire na948_9;
wire na949_1;
wire na950_1;
wire na950_2;
wire na951_2;
wire na952_2;
wire na953_1;
wire na953_9;
wire na954_2;
wire na955_1;
wire na955_2;
wire na956_1;
wire na957_2;
wire na958_1;
wire na959_2;
wire na960_1;
wire na960_2;
wire na961_1;
wire na962_2;
wire na963_1;
wire na963_2;
wire na964_2;
wire na965_1;
wire na966_1;
wire na967_2;
wire na968_1;
wire na968_2;
wire na969_1;
wire na970_1;
wire na971_1;
wire na972_2;
wire na973_1;
wire na973_2;
wire na974_2;
wire na975_1;
wire na976_1;
wire na977_2;
wire na978_1;
wire na979_2;
wire na980_1;
wire na980_2;
wire na981_1;
wire na982_1;
wire na982_2;
wire na983_2;
wire na984_2;
wire na985_2;
wire na986_1;
wire na987_1;
wire na987_2;
wire na988_1;
wire na989_2;
wire na990_2;
wire na991_1;
wire na992_2;
wire na993_1;
wire na995_1;
wire na995_2;
wire na996_1;
wire na998_2;
wire na1000_1;
wire na1000_2;
wire na1001_1;
wire na1003_2;
wire na1009_1;
wire na1010_1;
wire na1010_2;
wire na1011_2;
wire na1014_1;
wire na1015_1;
wire na1015_2;
wire na1016_2;
wire na1019_2;
wire na1020_1;
wire na1020_2;
wire na1021_1;
wire na1024_1;
wire na1025_1;
wire na1025_2;
wire na1026_1;
wire na1029_2;
wire na1030_1;
wire na1030_2;
wire na1031_1;
wire na1033_1;
wire na1033_2;
wire na1034_2;
wire na1036_1;
wire na1038_1;
wire na1038_2;
wire na1039_2;
wire na1041_1;
wire na1044_2;
wire na1045_1;
wire na1045_2;
wire na1046_1;
wire na1048_1;
wire na1048_2;
wire na1049_2;
wire na1051_1;
wire na1054_2;
wire na1055_1;
wire na1055_2;
wire na1056_2;
wire na1058_1;
wire na1059_2;
wire na1060_1;
wire na1060_2;
wire na1063_1;
wire na1063_2;
wire na1064_1;
wire na1066_2;
wire na1069_1;
wire na1070_1;
wire na1070_2;
wire na1071_1;
wire na1073_1;
wire na1073_2;
wire na1074_2;
wire na1076_1;
wire na1078_1;
wire na1078_2;
wire na1079_2;
wire na1081_1;
wire na1083_1;
wire na1083_2;
wire na1084_2;
wire na1086_1;
wire na1088_1;
wire na1088_2;
wire na1089_2;
wire na1091_2;
wire na1098_1;
wire na1098_2;
wire na1100_2;
wire na1101_1;
wire na1103_1;
wire na1103_2;
wire na1104_2;
wire na1106_1;
wire na1109_2;
wire na1110_1;
wire na1110_2;
wire na1111_1;
wire na1114_2;
wire na1115_1;
wire na1115_2;
wire na1116_1;
wire na1119_2;
wire na1120_1;
wire na1120_2;
wire na1121_1;
wire na1122_1;
wire na1122_2;
wire na1124_2;
wire na1125_1;
wire na1126_1;
wire na1126_2;
wire na1130_2;
wire na1131_1;
wire na1131_2;
wire na1132_1;
wire na1134_1;
wire na1134_2;
wire na1135_2;
wire na1137_1;
wire na1140_1;
wire na1141_1;
wire na1141_2;
wire na1142_1;
wire na1144_1;
wire na1144_2;
wire na1145_2;
wire na1147_1;
wire na1150_2;
wire na1151_1;
wire na1151_2;
wire na1152_1;
wire na1152_2;
wire na1156_1;
wire na1157_1;
wire na1157_2;
wire na1158_2;
wire na1160_1;
wire na1160_2;
wire na1161_1;
wire na1163_2;
wire na1165_1;
wire na1165_2;
wire na1166_2;
wire na1168_1;
wire na1175_2;
wire na1196_1;
wire na1198_2;
wire na1200_1;
wire na1201_2;
wire na1203_2;
wire na1204_2;
wire na1205_2;
wire na1206_2;
wire na1207_2;
wire na1208_2;
wire na1209_2;
wire na1210_2;
wire na1211_2;
wire na1212_2;
wire na1213_2;
wire na1214_2;
wire na1215_2;
wire na1216_2;
wire na1217_2;
wire na1218_2;
wire na1219_2;
wire na1220_2;
wire na1221_2;
wire na1222_2;
wire na1223_2;
wire na1224_2;
wire na1225_2;
wire na1226_2;
wire na1227_2;
wire na1228_2;
wire na1229_2;
wire na1230_2;
wire na1231_2;
wire na1232_2;
wire na1233_2;
wire na1234_2;
wire na1235_2;
wire na1236_2;
wire na1237_2;
wire na1238_2;
wire na1239_2;
wire na1240_2;
wire na1241_2;
wire na1242_2;
wire na1243_2;
wire na1244_2;
wire na1245_2;
wire na1246_2;
wire na1247_2;
wire na1248_2;
wire na1249_2;
wire na1250_2;
wire na1251_2;
wire na1252_2;
wire na1253_2;
wire na1254_2;
wire na1255_2;
wire na1256_2;
wire na1257_2;
wire na1258_2;
wire na1259_2;
wire na1260_2;
wire na1261_2;
wire na1262_2;
wire na1263_2;
wire na1264_2;
wire na1265_2;
wire na1266_2;
wire na1267_2;
wire na1268_2;
wire na1269_2;
wire na1270_2;
wire na1271_2;
wire na1272_2;
wire na1273_2;
wire na1274_2;
wire na1275_2;
wire na1276_2;
wire na1277_2;
wire na1278_2;
wire na1279_2;
wire na1280_2;
wire na1281_2;
wire na1282_2;
wire na879_25;
wire na879_26;
wire na879_27;
wire na879_28;
wire na879_29;
wire na879_30;
wire na879_31;
wire na879_32;
wire na879_33;
wire na879_34;
wire na879_35;
wire na879_36;
wire na879_37;
wire na879_38;
wire na879_39;
wire na879_40;
wire na908_10;
wire na910_10;
wire na915_10;
wire na918_10;
wire na923_10;
wire na929_10;
wire na934_10;
wire na937_10;
wire na947_10;
wire na952_10;
wire clk_check;
wire na1204_10;
wire na1205_10;
wire na1206_10;
wire na1207_10;
wire na1208_10;
wire na1209_10;
wire na1210_10;
wire na1211_10;
wire na1212_10;
wire na1213_10;
wire na1214_10;
wire na1215_10;
wire uart_rx_serial;

// C_ORAND*/D///      x90y45     80'h00_FA00_00_0000_0788_FD5D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1_1 ( .OUT(na1_1_i), .IN1(~na10_1), .IN2(na1216_2), .IN3(~na1217_2), .IN4(1'b0), .IN5(~na10_2), .IN6(na1216_2), .IN7(1'b1),
                   .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1_2 ( .OUT(na1_1), .CLK(na685_1), .EN(na270_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1_1_i) );
// C_AND///AND/      x89y49     80'h00_0078_00_0000_0C88_84AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3_1 ( .OUT(na3_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1268_2), .IN6(na7_2), .IN7(na4_2), .IN8(na704_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3_4 ( .OUT(na3_2), .IN1(na648_1), .IN2(1'b1), .IN3(na1220_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y43     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4_4 ( .OUT(na4_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na703_2), .IN4(na704_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x89y42     80'h00_0078_00_0000_0C88_8381
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a7_1 ( .OUT(na7_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na710_1), .IN7(na708_1), .IN8(na709_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7_4 ( .OUT(na7_2), .IN1(~na707_2), .IN2(~na710_1), .IN3(na708_1), .IN4(na709_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x90y43     80'h00_0078_00_0000_0C88_158F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1268_2), .IN6(1'b1), .IN7(~na703_2), .IN8(~na704_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8_4 ( .OUT(na8_2), .IN1(1'b1), .IN2(1'b1), .IN3(na703_2), .IN4(na704_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y43     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9_4 ( .OUT(na9_2), .IN1(na707_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na704_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x89y51     80'h00_0078_00_0000_0C88_88A8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a10_1 ( .OUT(na10_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1268_2), .IN6(na7_2), .IN7(na8_2), .IN8(na704_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a10_4 ( .OUT(na10_2), .IN1(na9_2), .IN2(na7_1), .IN3(na8_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x89y41     80'h00_FA00_00_0000_0EEE_A7AA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1_i), .IN1(na1225_2), .IN2(1'b0), .IN3(na900_1), .IN4(1'b0), .IN5(~na899_1), .IN6(~na17_1), .IN7(na13_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a12_2 ( .OUT(na12_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na12_1_i) );
// C_AND///AND/      x92y41     80'h00_0078_00_0000_0C88_F4F4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na12_1), .IN6(na22_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a13_4 ( .OUT(na13_2), .IN1(~na12_1), .IN2(na22_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y45     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a15_1 ( .OUT(na15_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na703_1), .IN8(~na704_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y48     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a17_1 ( .OUT(na17_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na18_1), .IN6(~na1152_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y47     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a18_1 ( .OUT(na18_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1268_2), .IN6(na7_2), .IN7(na4_2), .IN8(na704_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x89y50     80'h00_0078_00_0000_0C88_84A8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1268_2), .IN6(na7_2), .IN7(na8_2), .IN8(na704_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a22_4 ( .OUT(na22_2), .IN1(na15_1), .IN2(na7_2), .IN3(na8_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x92y40     80'h00_FA00_00_0000_0EEE_3C3E
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a23_1 ( .OUT(na23_1_i), .IN1(na903_2), .IN2(na905_2), .IN3(1'b0), .IN4(~na902_1), .IN5(1'b0), .IN6(na1152_2), .IN7(1'b0),
                    .IN8(~na902_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a23_2 ( .OUT(na23_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na23_1_i) );
// C_ORAND*/D///      x89y39     80'h00_FA00_00_0000_0788_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a27_1 ( .OUT(na27_1_i), .IN1(~na10_1), .IN2(~na651_1), .IN3(~na566_2), .IN4(~na1228_2), .IN5(~na10_2), .IN6(~na1252_2),
                    .IN7(~na343_2), .IN8(~na1230_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a27_2 ( .OUT(na27_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na27_1_i) );
// C_ORAND*/D///      x92y39     80'h00_FA00_00_0000_0788_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a30_1 ( .OUT(na30_1_i), .IN1(~na10_1), .IN2(~na651_2), .IN3(~na1227_2), .IN4(~na588_1), .IN5(~na10_2), .IN6(~na1253_2),
                    .IN7(~na1229_2), .IN8(~na365_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a30_2 ( .OUT(na30_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na30_1_i) );
// C_OR/D///      x89y37     80'h00_FA00_00_0000_0EEE_AD0D
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_1 ( .OUT(na33_1_i), .IN1(~na913_1), .IN2(na916_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na913_2), .IN6(na1152_2), .IN7(na914_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a33_2 ( .OUT(na33_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na33_1_i) );
// C_OR/D///      x82y35     80'h00_FA00_00_0000_0EEE_33DA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1_i), .IN1(na921_1), .IN2(1'b0), .IN3(~na37_2), .IN4(na919_1), .IN5(1'b0), .IN6(~na1270_2), .IN7(1'b0),
                    .IN8(~na920_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a36_2 ( .OUT(na36_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na36_1_i) );
// C_///AND/      x90y39     80'h00_0060_00_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a37_4 ( .OUT(na37_2), .IN1(~na18_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na43_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x83y39     80'h00_FA00_00_0000_0EEE_CB07
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a41_1 ( .OUT(na41_1_i), .IN1(~na42_2), .IN2(~na925_1), .IN3(1'b0), .IN4(1'b0), .IN5(na924_2), .IN6(~na925_2), .IN7(1'b0),
                    .IN8(na926_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a41_2 ( .OUT(na41_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na41_1_i) );
// C_///AND/      x89y47     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a42_4 ( .OUT(na42_2), .IN1(1'b1), .IN2(~na1152_2), .IN3(1'b1), .IN4(~na43_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x92y52     80'h00_0078_00_0000_0C88_8C8C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a43_1 ( .OUT(na43_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na7_2), .IN7(na4_2), .IN8(na704_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a43_4 ( .OUT(na43_2), .IN1(1'b1), .IN2(na7_2), .IN3(na8_1), .IN4(na704_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x83y42     80'h00_FA00_00_0000_0EEE_5ECC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a46_1 ( .OUT(na46_1_i), .IN1(1'b0), .IN2(na927_1), .IN3(1'b0), .IN4(na48_1), .IN5(na49_2), .IN6(na927_2), .IN7(~na37_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a46_2 ( .OUT(na46_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na46_1_i) );
// C_AND////      x94y40     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a48_1 ( .OUT(na48_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_1), .IN6(na7_2), .IN7(na8_2), .IN8(na392_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x83y41     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a49_4 ( .OUT(na49_2), .IN1(na9_2), .IN2(na7_1), .IN3(na8_1), .IN4(na456_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x90y37     80'h00_FA00_00_0000_0EEE_CDC5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a50_1 ( .OUT(na50_1_i), .IN1(~na930_1), .IN2(1'b0), .IN3(1'b0), .IN4(na53_1), .IN5(~na930_2), .IN6(na933_2), .IN7(1'b0),
                    .IN8(na931_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a50_2 ( .OUT(na50_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na50_1_i) );
// C_AND////      x92y44     80'h00_0018_00_0000_0C88_44FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a53_1 ( .OUT(na53_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1268_2), .IN6(na7_2), .IN7(~na703_2), .IN8(na704_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x90y36     80'h00_FA00_00_0000_0EEE_A70B
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a54_1 ( .OUT(na54_1_i), .IN1(na936_1), .IN2(~na938_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na56_1), .IN6(~na938_2), .IN7(na939_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a54_2 ( .OUT(na54_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na54_1_i) );
// C_AND////      x91y45     80'h00_0018_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a56_1 ( .OUT(na56_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na57_1), .IN8(~na43_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x94y47     80'h00_0018_00_0000_0888_536C
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a57_1 ( .OUT(na57_1), .IN1(1'b0), .IN2(~na7_2), .IN3(~na703_1), .IN4(na704_1), .IN5(1'b0), .IN6(na1269_2), .IN7(na703_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x83y44     80'h00_FA00_00_0000_0EEE_5E5A
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a59_1 ( .OUT(na59_1_i), .IN1(na3_1), .IN2(1'b0), .IN3(~na941_2), .IN4(1'b0), .IN5(na944_2), .IN6(na942_1), .IN7(~na941_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a59_2 ( .OUT(na59_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na59_1_i) );
// C_OR/D///      x80y43     80'h00_FA00_00_0000_0EEE_C0EB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a62_1 ( .OUT(na62_1_i), .IN1(na65_1), .IN2(~na17_1), .IN3(na64_2), .IN4(na945_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na945_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a62_2 ( .OUT(na62_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na62_1_i) );
// C_///AND/      x92y45     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a64_4 ( .OUT(na64_2), .IN1(na15_1), .IN2(na7_2), .IN3(na8_2), .IN4(na334_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y41     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a65_1 ( .OUT(na65_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9_2), .IN6(na7_1), .IN7(na8_1), .IN8(na397_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x81y37     80'h00_FA00_00_0000_0EEE_7AB0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a66_1 ( .OUT(na66_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na949_1), .IN4(~na950_1), .IN5(na951_2), .IN6(1'b0), .IN7(~na37_2),
                    .IN8(~na950_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a66_2 ( .OUT(na66_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na66_1_i) );
// C_OR/D///      x94y39     80'h00_FA00_00_0000_0EEE_555E
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a69_1 ( .OUT(na69_1_i), .IN1(na956_1), .IN2(na954_2), .IN3(~na955_1), .IN4(1'b0), .IN5(~na42_2), .IN6(1'b0), .IN7(~na955_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a69_2 ( .OUT(na69_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na69_1_i) );
// C_OR/D///      x83y47     80'h00_FA00_00_0000_0EEE_53E3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a72_1 ( .OUT(na72_1_i), .IN1(1'b0), .IN2(~na960_1), .IN3(na961_1), .IN4(na959_2), .IN5(1'b0), .IN6(~na960_2), .IN7(~na37_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a72_2 ( .OUT(na72_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na72_1_i) );
// C_OR/D///      x80y35     80'h00_FA00_00_0000_0EEE_E5A5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1_i), .IN1(~na963_1), .IN2(1'b0), .IN3(na966_1), .IN4(1'b0), .IN5(~na963_2), .IN6(1'b0), .IN7(na964_2),
                    .IN8(na53_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a75_2 ( .OUT(na75_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na75_1_i) );
// C_OR/D///      x81y40     80'h00_FA00_00_0000_0EEE_3E3A
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1_i), .IN1(na3_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na968_1), .IN5(na971_1), .IN6(na969_1), .IN7(1'b0), .IN8(~na968_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a78_2 ( .OUT(na78_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_1_i) );
// C_OR/D///      x90y41     80'h00_FA00_00_0000_0EEE_B0BA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a81_1 ( .OUT(na81_1_i), .IN1(na974_2), .IN2(1'b0), .IN3(na976_1), .IN4(~na973_1), .IN5(1'b0), .IN6(1'b0), .IN7(na57_1),
                    .IN8(~na973_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a81_2 ( .OUT(na81_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na81_1_i) );
// C_OR/D///      x90y42     80'h00_FA00_00_0000_0EEE_53E5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a84_1 ( .OUT(na84_1_i), .IN1(~na56_1), .IN2(1'b0), .IN3(na981_1), .IN4(na979_2), .IN5(1'b0), .IN6(~na1276_2), .IN7(~na980_1),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a84_2 ( .OUT(na84_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na84_1_i) );
// C_OR/D///      x82y42     80'h00_FA00_00_0000_0EEE_C3EE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a87_1 ( .OUT(na87_1_i), .IN1(na3_1), .IN2(na985_2), .IN3(na1281_2), .IN4(na982_2), .IN5(1'b0), .IN6(~na984_2), .IN7(1'b0),
                    .IN8(na982_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a87_2 ( .OUT(na87_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na87_1_i) );
// C_OR/D///      x90y44     80'h00_FA00_00_0000_0EEE_D0DA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1_i), .IN1(na18_1), .IN2(1'b0), .IN3(~na987_2), .IN4(na990_2), .IN5(1'b0), .IN6(1'b0), .IN7(~na987_1),
                    .IN8(na988_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a90_2 ( .OUT(na90_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na90_1_i) );
// C_ORAND*/D///      x83y49     80'h00_FA00_00_0000_0788_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a93_1 ( .OUT(na93_1_i), .IN1(~na1258_2), .IN2(~na22_1), .IN3(~na345_1), .IN4(~na1230_2), .IN5(~na10_1), .IN6(~na1264_2),
                    .IN7(~na408_2), .IN8(~na1224_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a93_2 ( .OUT(na93_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na93_1_i) );
// C_OR/D///      x90y47     80'h00_FA00_00_0000_0EEE_3C3E
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a96_1 ( .OUT(na96_1_i), .IN1(na996_1), .IN2(na998_2), .IN3(1'b0), .IN4(~na995_2), .IN5(1'b0), .IN6(na1152_2), .IN7(1'b0),
                    .IN8(~na995_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a96_2 ( .OUT(na96_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na96_1_i) );
// C_OR/D///      x83y43     80'h00_FA00_00_0000_0EEE_DCD0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a99_1 ( .OUT(na99_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1000_1), .IN4(na1003_2), .IN5(1'b0), .IN6(na1152_2), .IN7(~na1000_2),
                    .IN8(na1001_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a99_2 ( .OUT(na99_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na99_1_i) );
// C_ORAND*/D///      x83y45     80'h00_FA00_00_0000_0788_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a102_1 ( .OUT(na102_1_i), .IN1(~na1259_2), .IN2(~na22_1), .IN3(~na412_1), .IN4(~na1224_2), .IN5(~na10_1), .IN6(~na1265_2),
                     .IN7(~na1229_2), .IN8(~na347_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a102_2 ( .OUT(na102_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na102_1_i) );
// C_OR/D///      x82y48     80'h00_FA00_00_0000_0EEE_DC55
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a105_1 ( .OUT(na105_1_i), .IN1(~na107_2), .IN2(1'b0), .IN3(~na1010_2), .IN4(1'b0), .IN5(1'b0), .IN6(na1009_1), .IN7(~na1010_1),
                     .IN8(na1011_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a105_2 ( .OUT(na105_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na105_1_i) );
// C_///AND/      x89y53     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a107_4 ( .OUT(na107_2), .IN1(~na18_1), .IN2(1'b1), .IN3(~na57_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x83y48     80'h00_FA00_00_0000_0EEE_DC55
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a109_1 ( .OUT(na109_1_i), .IN1(~na42_2), .IN2(1'b0), .IN3(~na1015_2), .IN4(1'b0), .IN5(1'b0), .IN6(na1016_2), .IN7(~na1015_1),
                     .IN8(na1014_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a109_2 ( .OUT(na109_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na109_1_i) );
// C_OR/D///      x82y49     80'h00_FA00_00_0000_0EEE_C5C7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a112_1 ( .OUT(na112_1_i), .IN1(~na1020_1), .IN2(~na1236_2), .IN3(1'b0), .IN4(na1019_2), .IN5(~na1020_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na1021_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a112_2 ( .OUT(na112_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na112_1_i) );
// C_OR/D///      x83y50     80'h00_FA00_00_0000_0EEE_DA55
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a115_1 ( .OUT(na115_1_i), .IN1(~na117_1), .IN2(1'b0), .IN3(~na1025_2), .IN4(1'b0), .IN5(na1024_1), .IN6(1'b0), .IN7(~na1025_1),
                     .IN8(na1026_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a115_2 ( .OUT(na115_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na115_1_i) );
// C_AND////      x91y49     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a117_1 ( .OUT(na117_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3_1), .IN6(1'b1), .IN7(~na57_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x90y49     80'h00_FA00_00_0000_0EEE_CD33
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a119_1 ( .OUT(na119_1_i), .IN1(1'b0), .IN2(~na1280_2), .IN3(1'b0), .IN4(~na1030_2), .IN5(~na56_1), .IN6(na1029_2), .IN7(1'b0),
                     .IN8(na1031_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a119_2 ( .OUT(na119_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na119_1_i) );
// C_OR/D///      x83y52     80'h00_FA00_00_0000_0EEE_BC3A
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a122_1 ( .OUT(na122_1_i), .IN1(na3_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1033_2), .IN5(1'b0), .IN6(na1034_2), .IN7(na1036_1),
                     .IN8(~na1033_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a122_2 ( .OUT(na122_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na122_1_i) );
// C_OR/D///      x90y52     80'h00_FA00_00_0000_0EEE_30BE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a125_1 ( .OUT(na125_1_i), .IN1(na18_1), .IN2(na1039_2), .IN3(na1041_1), .IN4(~na1038_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(~na1038_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a125_2 ( .OUT(na125_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na125_1_i) );
// C_OR/D///      x83y51     80'h00_FA00_00_0000_0EEE_A5D5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1_i), .IN1(~na1045_2), .IN2(1'b0), .IN3(~na37_2), .IN4(na1044_2), .IN5(~na1045_1), .IN6(1'b0), .IN7(na1046_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a128_2 ( .OUT(na128_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na128_1_i) );
// C_OR/D///      x90y53     80'h00_FA00_00_0000_0EEE_C5E5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a131_1 ( .OUT(na131_1_i), .IN1(~na1048_1), .IN2(1'b0), .IN3(na1051_1), .IN4(na1049_2), .IN5(~na1048_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na43_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a131_2 ( .OUT(na131_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na131_1_i) );
// C_OR/D///      x83y53     80'h00_FA00_00_0000_0EEE_C7C3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a134_1 ( .OUT(na134_1_i), .IN1(1'b0), .IN2(~na1055_1), .IN3(1'b0), .IN4(na1054_2), .IN5(~na107_2), .IN6(~na1055_2), .IN7(1'b0),
                     .IN8(na1056_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a134_2 ( .OUT(na134_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na134_1_i) );
// C_OR/D///      x80y51     80'h00_FA00_00_0000_0EEE_CDC3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a137_1 ( .OUT(na137_1_i), .IN1(1'b0), .IN2(~na1058_1), .IN3(1'b0), .IN4(na138_2), .IN5(~na117_1), .IN6(na1059_2), .IN7(1'b0),
                     .IN8(na138_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a137_2 ( .OUT(na137_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na137_1_i) );
// C_AND///AND/      x90y48     80'h00_0078_00_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(1'b1), .IN8(na360_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a138_4 ( .OUT(na138_2), .IN1(1'b1), .IN2(na22_1), .IN3(1'b1), .IN4(na583_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x89y54     80'h00_FA00_00_0000_0EEE_CEAE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a141_1 ( .OUT(na141_1_i), .IN1(na3_1), .IN2(na1060_1), .IN3(na1281_2), .IN4(1'b0), .IN5(na3_2), .IN6(na1060_2), .IN7(1'b0),
                     .IN8(na145_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a141_2 ( .OUT(na141_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na141_1_i) );
// C_///AND/      x90y50     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a145_4 ( .OUT(na145_2), .IN1(na15_1), .IN2(na7_2), .IN3(na8_2), .IN4(na360_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x90y54     80'h00_FA00_00_0000_0EEE_ABA3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a146_1 ( .OUT(na146_1_i), .IN1(1'b0), .IN2(~na1063_1), .IN3(na1066_2), .IN4(1'b0), .IN5(na1064_1), .IN6(~na1063_2), .IN7(na57_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a146_2 ( .OUT(na146_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na146_1_i) );
// C_OR/D///      x83y55     80'h00_FA00_00_0000_0EEE_C5A7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a149_1 ( .OUT(na149_1_i), .IN1(~na1070_1), .IN2(~na1233_2), .IN3(na1069_1), .IN4(1'b0), .IN5(~na1070_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na1071_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a149_2 ( .OUT(na149_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na149_1_i) );
// C_OR/D///      x94y57     80'h00_FA00_00_0000_0EEE_BAB0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a152_1 ( .OUT(na152_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1076_1), .IN4(~na1073_2), .IN5(na3_1), .IN6(1'b0), .IN7(na1074_2),
                     .IN8(~na1073_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a152_2 ( .OUT(na152_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na152_1_i) );
// C_OR/D///      x89y56     80'h00_FA00_00_0000_0EEE_BC3A
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a155_1 ( .OUT(na155_1_i), .IN1(na18_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1078_2), .IN5(1'b0), .IN6(na1079_2), .IN7(na1081_1),
                     .IN8(~na1078_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a155_2 ( .OUT(na155_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na155_1_i) );
// C_OR/D///      x90y56     80'h00_FA00_00_0000_0EEE_0BE3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a158_1 ( .OUT(na158_1_i), .IN1(1'b0), .IN2(~na1083_1), .IN3(na1281_2), .IN4(na1086_1), .IN5(na1084_2), .IN6(~na1083_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a158_2 ( .OUT(na158_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na158_1_i) );
// C_OR/D///      x83y57     80'h00_FA00_00_0000_0EEE_DC5C
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a161_1 ( .OUT(na161_1_i), .IN1(1'b0), .IN2(na1091_2), .IN3(~na1088_2), .IN4(1'b0), .IN5(1'b0), .IN6(na1152_2), .IN7(~na1088_1),
                     .IN8(na1089_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a161_2 ( .OUT(na161_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na161_1_i) );
// C_ORAND*/D///      x89y57     80'h00_FA00_00_0000_0788_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a164_1 ( .OUT(na164_1_i), .IN1(~na1260_2), .IN2(~na22_1), .IN3(~na1229_2), .IN4(~na369_1), .IN5(~na10_1), .IN6(~na655_2),
                     .IN7(~na1223_2), .IN8(~na432_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a164_2 ( .OUT(na164_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na164_1_i) );
// C_ORAND*/D///      x90y57     80'h00_FA00_00_0000_0788_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a167_1 ( .OUT(na167_1_i), .IN1(~na1261_2), .IN2(~na22_1), .IN3(~na434_1), .IN4(~na1224_2), .IN5(~na10_1), .IN6(~na1266_2),
                     .IN7(~na1229_2), .IN8(~na369_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a167_2 ( .OUT(na167_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na167_1_i) );
// C_OR/D///      x83y58     80'h00_FA00_00_0000_0EEE_3CEE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a170_1 ( .OUT(na170_1_i), .IN1(na18_1), .IN2(na1098_1), .IN3(na1101_1), .IN4(na43_2), .IN5(1'b0), .IN6(na1098_2), .IN7(1'b0),
                     .IN8(~na1100_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a170_2 ( .OUT(na170_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na170_1_i) );
// C_OR/D///      x89y58     80'h00_FA00_00_0000_0EEE_E3C3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a173_1 ( .OUT(na173_1_i), .IN1(1'b0), .IN2(~na1103_1), .IN3(1'b0), .IN4(na43_1), .IN5(1'b0), .IN6(~na1103_2), .IN7(na1104_2),
                     .IN8(na1106_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a173_2 ( .OUT(na173_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na173_1_i) );
// C_OR/D///      x90y58     80'h00_FA00_00_0000_0EEE_3DB0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a176_1 ( .OUT(na176_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1109_2), .IN4(~na1110_2), .IN5(~na107_2), .IN6(na1111_1), .IN7(1'b0),
                     .IN8(~na1110_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a176_2 ( .OUT(na176_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na176_1_i) );
// C_OR/D///      x83y59     80'h00_FA00_00_0000_0EEE_BC35
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a179_1 ( .OUT(na179_1_i), .IN1(~na117_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1115_2), .IN5(1'b0), .IN6(na1116_1), .IN7(na1114_2),
                     .IN8(~na1115_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a179_2 ( .OUT(na179_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na179_1_i) );
// C_OR/D///      x89y59     80'h00_FA00_00_0000_0EEE_C5ED
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_1 ( .OUT(na182_1_i), .IN1(~na1120_1), .IN2(na1231_2), .IN3(na1119_2), .IN4(na43_2), .IN5(~na1120_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na1121_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a182_2 ( .OUT(na182_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na182_1_i) );
// C_OR/D///      x90y59     80'h00_FA00_00_0000_0EEE_ABCE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a186_1 ( .OUT(na186_1_i), .IN1(na1122_2), .IN2(na1152_2), .IN3(1'b0), .IN4(na1125_1), .IN5(na1122_1), .IN6(~na1124_2), .IN7(na1217_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a186_2 ( .OUT(na186_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na186_1_i) );
// C_OR/D///      x91y57     80'h00_FA00_00_0000_0EEE_E3AA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a189_1 ( .OUT(na189_1_i), .IN1(na191_1), .IN2(1'b0), .IN3(na1126_2), .IN4(1'b0), .IN5(1'b0), .IN6(~na17_1), .IN7(na1126_1),
                     .IN8(na192_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a189_2 ( .OUT(na189_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na189_1_i) );
// C_AND////      x93y49     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a191_1 ( .OUT(na191_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na15_1), .IN6(na7_2), .IN7(na8_2), .IN8(na378_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y50     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a192_4 ( .OUT(na192_2), .IN1(na9_2), .IN2(na7_1), .IN3(na8_1), .IN4(na441_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x89y60     80'h00_FA00_00_0000_0EEE_07AB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a193_1 ( .OUT(na193_1_i), .IN1(na1130_2), .IN2(~na1131_2), .IN3(na1132_1), .IN4(1'b0), .IN5(~na107_2), .IN6(~na1131_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a193_2 ( .OUT(na193_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na193_1_i) );
// C_OR/D///      x90y60     80'h00_FA00_00_0000_0EEE_DCD0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a196_1 ( .OUT(na196_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1134_1), .IN4(na1137_1), .IN5(1'b0), .IN6(na1231_2), .IN7(~na1134_2),
                     .IN8(na1135_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a196_2 ( .OUT(na196_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na196_1_i) );
// C_OR/D///      x81y63     80'h00_FA00_00_0000_0EEE_35BA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a199_1 ( .OUT(na199_1_i), .IN1(na1142_1), .IN2(1'b0), .IN3(na1140_1), .IN4(~na1141_2), .IN5(~na107_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(~na1141_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a199_2 ( .OUT(na199_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na199_1_i) );
// C_OR/D///      x89y61     80'h00_FA00_00_0000_0EEE_C5CD
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a202_1 ( .OUT(na202_1_i), .IN1(~na1144_2), .IN2(na1147_1), .IN3(1'b0), .IN4(na53_1), .IN5(~na1144_1), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na1145_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a202_2 ( .OUT(na202_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na202_1_i) );
// C_OR/D///      x90y61     80'h00_FA00_00_0000_0EEE_5EDC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a205_1 ( .OUT(na205_1_i), .IN1(1'b0), .IN2(na1152_1), .IN3(~na1151_1), .IN4(na1150_2), .IN5(na3_1), .IN6(na1152_2), .IN7(~na1151_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a205_2 ( .OUT(na205_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na205_1_i) );
// C_OR/D///      x91y60     80'h00_FA00_00_0000_0EEE_CBE3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a209_1 ( .OUT(na209_1_i), .IN1(1'b0), .IN2(~na1157_1), .IN3(na1156_1), .IN4(na43_2), .IN5(na1158_2), .IN6(~na1157_2), .IN7(1'b0),
                     .IN8(na43_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a209_2 ( .OUT(na209_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na209_1_i) );
// C_OR/D///      x82y61     80'h00_FA00_00_0000_0EEE_DAD0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a212_1 ( .OUT(na212_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na1160_2), .IN4(na1163_2), .IN5(na3_1), .IN6(1'b0), .IN7(~na1160_1),
                     .IN8(na1161_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a212_2 ( .OUT(na212_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na212_1_i) );
// C_OR/D///      x89y62     80'h00_FA00_00_0000_0EEE_07CE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a215_1 ( .OUT(na215_1_i), .IN1(na1168_1), .IN2(na1166_2), .IN3(1'b0), .IN4(na1226_2), .IN5(~na1282_2), .IN6(~na1165_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a215_2 ( .OUT(na215_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na215_1_i) );
// C_ORAND*/D///      x80y59     80'h00_FA00_00_0000_0788_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a218_1 ( .OUT(na218_1_i), .IN1(~na1262_2), .IN2(~na22_1), .IN3(~na389_1), .IN4(~na1230_2), .IN5(~na10_1), .IN6(~na1267_2),
                     .IN7(~na452_2), .IN8(~na1224_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a218_2 ( .OUT(na218_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na218_1_i) );
// C_ORAND*/D///      x83y63     80'h00_FA00_00_0000_0788_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a221_1 ( .OUT(na221_1_i), .IN1(~na1263_2), .IN2(~na22_1), .IN3(~na1223_2), .IN4(~na454_1), .IN5(~na10_1), .IN6(~na677_1),
                     .IN7(~na389_2), .IN8(~na1230_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a221_2 ( .OUT(na221_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na221_1_i) );
// C_MX2b/D///      x79y66     80'h00_ED00_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a224_1 ( .OUT(na224_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na784_1), .IN5(1'b0), .IN6(na878_1), .IN7(1'b0), .IN8(na873_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a224_2 ( .OUT(na224_1), .CLK(~na685_3), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na224_1_i) );
// C_AND////      x94y38     80'h00_0018_00_0000_0888_14A4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a227_1 ( .OUT(na227_1), .IN1(~na247_1), .IN2(na230_2), .IN3(na231_1), .IN4(1'b1), .IN5(~na247_2), .IN6(na229_1), .IN7(~na249_2),
                     .IN8(~na250_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y32     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a229_1 ( .OUT(na229_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na239_2), .IN6(~na236_1), .IN7(~na1243_2),
                     .IN8(~na237_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x89y34     80'h00_0060_00_0000_0C08_FF41
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a230_4 ( .OUT(na230_2), .IN1(~na1246_2), .IN2(~na245_1), .IN3(~na246_2), .IN4(na243_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y33     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a231_1 ( .OUT(na231_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na239_1), .IN6(~na241_2), .IN7(na1244_2), .IN8(~na243_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y33     80'h00_0018_00_0000_0C88_1AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a232_1 ( .OUT(na232_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na251_1), .IN6(1'b1), .IN7(~na258_1), .IN8(~na260_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x91y34     80'h00_0078_00_0000_0C88_2413
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a233_1 ( .OUT(na233_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na234_1), .IN6(na901_1), .IN7(na258_1), .IN8(~na260_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a233_4 ( .OUT(na233_2), .IN1(1'b1), .IN2(~na257_1), .IN3(~na857_1), .IN4(~na260_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y37     80'h00_0018_00_0000_0888_14A4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a234_1 ( .OUT(na234_1), .IN1(~na247_1), .IN2(na229_1), .IN3(na235_2), .IN4(1'b1), .IN5(~na247_2), .IN6(na230_2), .IN7(~na249_2),
                     .IN8(~na250_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y29     80'h00_0060_00_0000_0C08_FF81
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a235_4 ( .OUT(na235_2), .IN1(~na239_1), .IN2(~na241_1), .IN3(na1245_2), .IN4(na243_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x89y28     80'h00_FA00_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a236_1 ( .OUT(na236_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1175_2), .IN6(1'b1), .IN7(na542_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a236_2 ( .OUT(na236_1), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na236_1_i) );
// C_AND/D//AND/D      x90y30     80'h00_FA00_80_0000_0C88_A535
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a237_1 ( .OUT(na237_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1175_2), .IN6(1'b1), .IN7(na542_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a237_2 ( .OUT(na237_1), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na237_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a237_4 ( .OUT(na237_2_i), .IN1(~na1175_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na237_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a237_5 ( .OUT(na237_2), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na237_2_i) );
// C_AND/D//AND/D      x91y33     80'h00_FA00_80_0000_0C88_C5C5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a239_1 ( .OUT(na239_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1175_2), .IN6(1'b1), .IN7(1'b1), .IN8(na544_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a239_2 ( .OUT(na239_1), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na239_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a239_4 ( .OUT(na239_2_i), .IN1(~na1175_2), .IN2(1'b1), .IN3(1'b1), .IN4(na544_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a239_5 ( .OUT(na239_2), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na239_2_i) );
// C_AND/D//AND/D      x87y32     80'h00_FA00_80_0000_0C88_A5A5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a241_1 ( .OUT(na241_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1175_2), .IN6(1'b1), .IN7(na546_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a241_2 ( .OUT(na241_1), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na241_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a241_4 ( .OUT(na241_2_i), .IN1(~na1175_2), .IN2(1'b1), .IN3(na546_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a241_5 ( .OUT(na241_2), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na241_2_i) );
// C_AND/D//AND/D      x90y32     80'h00_FA00_80_0000_0C88_C5C5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a243_1 ( .OUT(na243_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1175_2), .IN6(1'b1), .IN7(1'b1), .IN8(na548_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a243_2 ( .OUT(na243_1), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na243_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a243_4 ( .OUT(na243_2_i), .IN1(~na1175_2), .IN2(1'b1), .IN3(1'b1), .IN4(na548_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a243_5 ( .OUT(na243_2), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na243_2_i) );
// C_AND/D//AND/D      x91y30     80'h00_FA00_80_0000_0C88_A5A5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a245_1 ( .OUT(na245_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1175_2), .IN6(1'b1), .IN7(na550_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a245_2 ( .OUT(na245_1), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na245_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a245_4 ( .OUT(na245_2_i), .IN1(~na1175_2), .IN2(1'b1), .IN3(na550_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a245_5 ( .OUT(na245_2), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na245_2_i) );
// C_///AND/D      x94y35     80'h00_FA00_80_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a246_4 ( .OUT(na246_2_i), .IN1(~na1175_2), .IN2(1'b1), .IN3(1'b1), .IN4(na537_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a246_5 ( .OUT(na246_2), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na246_2_i) );
// C_AND/D//AND/D      x95y35     80'h00_FA00_80_0000_0C88_C5A5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a247_1 ( .OUT(na247_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1175_2), .IN6(1'b1), .IN7(1'b1), .IN8(na537_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a247_2 ( .OUT(na247_1), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na247_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a247_4 ( .OUT(na247_2_i), .IN1(~na1175_2), .IN2(1'b1), .IN3(na539_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a247_5 ( .OUT(na247_2), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na247_2_i) );
// C_///AND/D      x94y37     80'h00_FA00_80_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a249_4 ( .OUT(na249_2_i), .IN1(~na1175_2), .IN2(1'b1), .IN3(na539_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a249_5 ( .OUT(na249_2), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na249_2_i) );
// C_///AND/D      x94y34     80'h00_FA00_80_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a250_4 ( .OUT(na250_2_i), .IN1(~na1175_2), .IN2(1'b1), .IN3(1'b1), .IN4(na541_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a250_5 ( .OUT(na250_2), .CLK(na685_1), .EN(na266_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na250_2_i) );
// C_ORAND*/D///      x89y35     80'h00_FE00_00_0000_0788_D357
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a251_1 ( .OUT(na251_1_i), .IN1(~na251_1), .IN2(~na233_1), .IN3(~na252_1), .IN4(1'b0), .IN5(1'b0), .IN6(~na233_2), .IN7(~na1242_2),
                     .IN8(na227_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a251_2 ( .OUT(na251_1), .CLK(na685_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na251_1_i) );
// C_AND////      x86y33     80'h00_0018_00_0000_0888_F8C2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a252_1 ( .OUT(na252_1), .IN1(na265_2), .IN2(~na261_2), .IN3(1'b1), .IN4(na254_1), .IN5(na265_1), .IN6(na262_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x84y32     80'h00_0060_00_0000_0C08_FFC8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a253_4 ( .OUT(na253_2), .IN1(na265_1), .IN2(na262_1), .IN3(1'b1), .IN4(na1250_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y34     80'h00_0018_00_0000_0C88_25FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a254_1 ( .OUT(na254_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na251_1), .IN6(1'b1), .IN7(na258_1), .IN8(~na260_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*////D      x89y38     80'h00_FA18_00_0000_0788_F55F
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a257_1 ( .OUT(na257_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na258_1), .IN4(1'b1), .IN5(~na251_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a257_5 ( .OUT(na257_2), .CLK(na685_1), .EN(na268_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na257_1) );
// C_OR/D///      x90y33     80'h00_FE00_00_0000_0CEE_CE00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a258_1 ( .OUT(na258_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na259_1), .IN6(na233_1), .IN7(1'b0), .IN8(na254_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a258_2 ( .OUT(na258_1), .CLK(na685_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na258_1_i) );
// C_AND////      x89y31     80'h00_0018_00_0000_0C88_4AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a259_1 ( .OUT(na259_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na232_1), .IN6(1'b1), .IN7(~na857_1), .IN8(na227_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////D      x88y32     80'h00_FE18_00_0000_0888_F32A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a260_1 ( .OUT(na260_1), .IN1(na251_1), .IN2(1'b1), .IN3(na258_1), .IN4(~na260_2), .IN5(1'b1), .IN6(~na261_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a260_5 ( .OUT(na260_2), .CLK(na685_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na260_1) );
// C_///AND/      x89y36     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a261_4 ( .OUT(na261_2), .IN1(~na234_1), .IN2(na901_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x83y30     80'h00_F600_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a262_1 ( .OUT(na262_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na263_1), .IN7(na533_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a262_2 ( .OUT(na262_1), .CLK(na685_1), .EN(~na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na262_1_i) );
// C_AND////      x85y32     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a263_1 ( .OUT(na263_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1247_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na253_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x83y31     80'h00_F600_80_0000_0C88_ACF4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a265_1 ( .OUT(na265_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na263_1), .IN7(na533_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a265_2 ( .OUT(na265_1), .CLK(na685_1), .EN(~na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na265_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a265_4 ( .OUT(na265_2_i), .IN1(~na265_2), .IN2(na263_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a265_5 ( .OUT(na265_2), .CLK(na685_1), .EN(~na269_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na265_2_i) );
// C_///AND/      x94y33     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a266_4 ( .OUT(na266_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1196_1), .IN4(~na260_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x88y33     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a267_1 ( .OUT(na267_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na261_2), .IN7(1'b1), .IN8(na254_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x89y32     80'h00_0018_00_0040_0C24_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a268_1 ( .OUT(na268_1), .IN1(1'b0), .IN2(1'b1), .IN3(na1198_2), .IN4(1'b0), .IN5(~na251_1), .IN6(1'b1), .IN7(na258_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x86y32     80'h00_0018_00_0000_0C88_5EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a269_1 ( .OUT(na269_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1248_2), .IN6(na257_1), .IN7(~na267_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y45     80'h00_0060_00_0000_0C08_FF32
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a270_4 ( .OUT(na270_2), .IN1(na271_1), .IN2(~na22_2), .IN3(1'b1), .IN4(~na1228_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x91y53     80'h00_FE00_80_0000_0C88_F4FC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a271_1 ( .OUT(na271_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na271_2), .IN6(na257_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a271_2 ( .OUT(na271_1), .CLK(na685_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na271_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a271_4 ( .OUT(na271_2_i), .IN1(1'b1), .IN2(na257_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a271_5 ( .OUT(na271_2), .CLK(na685_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na271_2_i) );
// C_MX2b/D///      x85y33     80'h00_FA00_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a272_1 ( .OUT(na272_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na273_1), .IN4(1'b1), .IN5(na272_1), .IN6(1'b0), .IN7(na857_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a272_2 ( .OUT(na272_1), .CLK(na685_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na272_1_i) );
// C_AND////      x86y29     80'h00_0018_00_0000_0C88_21FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a273_1 ( .OUT(na273_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na265_2), .IN6(~na1257_2), .IN7(na912_1), .IN8(~na552_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x87y31     80'h00_FA00_00_0040_0C05_8000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a274_1 ( .OUT(na274_1_i), .IN1(na274_1), .IN2(1'b0), .IN3(na857_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na275_2), .IN8(na552_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a274_2 ( .OUT(na274_1), .CLK(na685_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na274_1_i) );
// C_///AND/      x86y31     80'h00_0060_00_0000_0C08_FF4A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a275_4 ( .OUT(na275_2), .IN1(na265_2), .IN2(1'b1), .IN3(~na912_1), .IN4(na552_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x91y35     80'h00_FA00_00_0040_0C05_8000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a276_1 ( .OUT(na276_1_i), .IN1(na276_1), .IN2(1'b0), .IN3(na857_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na277_1), .IN8(na552_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a276_2 ( .OUT(na276_1), .CLK(na685_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na276_1_i) );
// C_AND////      x86y31     80'h00_0018_00_0000_0C88_45FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a277_1 ( .OUT(na277_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na265_2), .IN6(1'b1), .IN7(~na912_1), .IN8(na552_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x91y29     80'h00_FA00_00_0040_0C05_8000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a278_1 ( .OUT(na278_1_i), .IN1(na278_1), .IN2(1'b0), .IN3(na857_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na279_2), .IN8(na552_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a278_2 ( .OUT(na278_1), .CLK(na685_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na278_1_i) );
// C_///AND/      x84y29     80'h00_0060_00_0000_0C08_FF1A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a279_4 ( .OUT(na279_2), .IN1(na265_2), .IN2(1'b1), .IN3(~na912_1), .IN4(~na552_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x85y29     80'h00_FA00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a280_1 ( .OUT(na280_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na281_2), .IN5(na280_1), .IN6(1'b0), .IN7(na857_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a280_2 ( .OUT(na280_1), .CLK(na685_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na280_1_i) );
// C_///AND/      x86y32     80'h00_0060_00_0000_0C08_FF14
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a281_4 ( .OUT(na281_2), .IN1(~na265_2), .IN2(na1257_2), .IN3(~na912_1), .IN4(~na552_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x87y27     80'h00_FA00_00_0040_0C05_2000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a282_1 ( .OUT(na282_1_i), .IN1(na282_1), .IN2(1'b0), .IN3(na857_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na275_2), .IN8(~na552_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a282_2 ( .OUT(na282_1), .CLK(na685_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na282_1_i) );
// C_MX2a/D///      x87y29     80'h00_FA00_00_0040_0C05_2000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a283_1 ( .OUT(na283_1_i), .IN1(na283_1), .IN2(1'b0), .IN3(na857_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na277_1), .IN8(~na552_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a283_2 ( .OUT(na283_1), .CLK(na685_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na283_1_i) );
// C_MX2a/D///      x83y29     80'h00_FA00_00_0040_0C05_2000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_1 ( .OUT(na284_1_i), .IN1(na284_1), .IN2(1'b0), .IN3(na857_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na279_2), .IN8(~na552_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_2 ( .OUT(na284_1), .CLK(na685_1), .EN(na267_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na284_1_i) );
// C_ORAND*/D///      x82y63     80'h00_FA00_00_0000_0788_F733
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a315_1 ( .OUT(na315_1_i), .IN1(1'b0), .IN2(~na1203_2), .IN3(1'b0), .IN4(~na43_2), .IN5(~na10_2), .IN6(~na1254_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a315_2 ( .OUT(na315_1), .CLK(na685_1), .EN(na271_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na315_1_i) );
// C_ADDF2///ADDF2/      x93y35     80'h00_0078_00_0020_0C66_5005
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a318_1 ( .OUT(na318_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na246_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na331_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a318_4 ( .OUT(na318_2), .COUTY1(na318_4), .IN1(~na247_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na246_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na331_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x93y36     80'h00_0078_00_0020_0C66_0550
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a320_1 ( .OUT(na320_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na247_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na318_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a320_4 ( .OUT(na320_2), .COUTY1(na320_4), .IN1(1'b0), .IN2(1'b0), .IN3(~na249_2), .IN4(1'b1), .IN5(~na247_2), .IN6(1'b1),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na318_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x93y37     80'h00_0018_00_0010_0666_0030
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a322_1 ( .OUT(na322_1), .COUTY1(na322_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na250_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na320_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x93y30     80'h00_0078_00_0020_0C66_3330
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a323_1 ( .OUT(na323_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na236_1), .IN7(1'b1), .IN8(~na237_2),
                     .CINX(1'b0), .CINY1(na332_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a323_4 ( .OUT(na323_2), .COUTY1(na323_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na237_1), .IN5(1'b1), .IN6(~na236_1),
                     .IN7(1'b1), .IN8(~na237_2), .CINX(1'b0), .CINY1(na332_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x93y31     80'h00_0078_00_0020_0C66_0505
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a325_1 ( .OUT(na325_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na239_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na323_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a325_4 ( .OUT(na325_2), .COUTY1(na325_4), .IN1(~na239_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na239_2), .IN6(1'b1),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na323_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x93y32     80'h00_0078_00_0020_0C66_F303
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a327_1 ( .OUT(na327_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na241_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na325_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a327_4 ( .OUT(na327_2), .COUTY1(na327_4), .IN1(1'b1), .IN2(~na241_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na241_2),
                     .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na325_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x93y33     80'h00_0078_00_0020_0C66_3F3F
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a329_1 ( .OUT(na329_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na243_2),
                     .CINX(1'b0), .CINY1(na327_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a329_4 ( .OUT(na329_2), .COUTY1(na329_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na243_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na243_2), .CINX(1'b0), .CINY1(na327_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x93y34     80'h00_0078_00_0020_0C66_0303
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a331_1 ( .OUT(na331_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na245_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na329_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a331_4 ( .OUT(na331_2), .COUTY1(na331_4), .IN1(1'b1), .IN2(~na245_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na245_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na329_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x93y29     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a332_2 ( .OUT(na332_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a332_6 ( .COUTY1(na332_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na332_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x84y38     80'h00_0078_00_0020_0C66_AF0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a334_1 ( .OUT(na334_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na62_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na394_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a334_4 ( .OUT(na334_2), .COUTY1(na334_4), .IN1(na66_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na62_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na394_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y39     80'h00_0078_00_0020_0C66_AF0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a336_1 ( .OUT(na336_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na69_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na334_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a336_4 ( .OUT(na336_2), .COUTY1(na336_4), .IN1(na72_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na69_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na334_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y40     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a338_1 ( .OUT(na338_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na75_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na336_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a338_4 ( .OUT(na338_2), .COUTY1(na338_4), .IN1(1'b1), .IN2(na78_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na75_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na336_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y41     80'h00_0078_00_0020_0C66_AFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a340_1 ( .OUT(na340_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na81_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na338_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a340_4 ( .OUT(na340_2), .COUTY1(na340_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na84_1), .IN5(1'b1), .IN6(1'b1), .IN7(na81_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na338_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y42     80'h00_0078_00_0020_0C66_CFC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a342_1 ( .OUT(na342_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                     .CINX(1'b0), .CINY1(na340_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a342_4 ( .OUT(na342_2), .COUTY1(na342_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na90_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na87_1), .CINX(1'b0), .CINY1(na340_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y33     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a343_1 ( .OUT(na343_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na12_1), .IN6(1'b1), .IN7(1'b1), .IN8(na23_1),
                     .CINX(1'b0), .CINY1(na395_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a343_4 ( .OUT(na343_2), .COUTY1(na343_4), .IN1(na27_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na12_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na23_1), .CINX(1'b0), .CINY1(na395_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y43     80'h00_0078_00_0020_0C66_0AAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a345_1 ( .OUT(na345_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na93_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na342_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a345_4 ( .OUT(na345_2), .COUTY1(na345_4), .IN1(1'b1), .IN2(1'b1), .IN3(na96_1), .IN4(1'b1), .IN5(na93_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na342_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y44     80'h00_0078_00_0020_0C66_FA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a347_1 ( .OUT(na347_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na99_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na345_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a347_4 ( .OUT(na347_2), .COUTY1(na347_4), .IN1(na102_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na99_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na345_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y45     80'h00_0078_00_0020_0C66_CFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a349_1 ( .OUT(na349_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na105_1),
                     .CINX(1'b0), .CINY1(na347_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a349_4 ( .OUT(na349_2), .COUTY1(na349_4), .IN1(1'b1), .IN2(na109_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na105_1), .CINX(1'b0), .CINY1(na347_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y46     80'h00_0078_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a351_1 ( .OUT(na351_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na112_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na349_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a351_4 ( .OUT(na351_2), .COUTY1(na351_4), .IN1(1'b1), .IN2(na115_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na112_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na349_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y47     80'h00_0078_00_0020_0C66_AF0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a353_1 ( .OUT(na353_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na119_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na351_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a353_4 ( .OUT(na353_2), .COUTY1(na353_4), .IN1(1'b1), .IN2(na122_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na119_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na351_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y48     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a356_1 ( .OUT(na356_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na125_1),
                     .CINX(1'b0), .CINY1(na353_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a356_4 ( .OUT(na356_2), .COUTY1(na356_4), .IN1(na128_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na125_1), .CINX(1'b0), .CINY1(na353_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y49     80'h00_0078_00_0020_0C66_A0FA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a358_1 ( .OUT(na358_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na131_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na356_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a358_4 ( .OUT(na358_2), .COUTY1(na358_4), .IN1(na134_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na131_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na356_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y50     80'h00_0078_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a360_1 ( .OUT(na360_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na137_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na358_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a360_4 ( .OUT(na360_2), .COUTY1(na360_4), .IN1(1'b1), .IN2(na141_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na137_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na358_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y51     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a362_1 ( .OUT(na362_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na146_1),
                     .CINX(1'b0), .CINY1(na360_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a362_4 ( .OUT(na362_2), .COUTY1(na362_4), .IN1(na149_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na146_1), .CINX(1'b0), .CINY1(na360_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y52     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a364_1 ( .OUT(na364_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na152_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na362_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a364_4 ( .OUT(na364_2), .COUTY1(na364_4), .IN1(1'b1), .IN2(na155_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na152_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na362_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y34     80'h00_0078_00_0020_0C66_A0FA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a365_1 ( .OUT(na365_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na30_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na343_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a365_4 ( .OUT(na365_2), .COUTY1(na365_4), .IN1(na33_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na30_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na343_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y53     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a367_1 ( .OUT(na367_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na158_1),
                     .CINX(1'b0), .CINY1(na364_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a367_4 ( .OUT(na367_2), .COUTY1(na367_4), .IN1(na161_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na158_1), .CINX(1'b0), .CINY1(na364_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y54     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a369_1 ( .OUT(na369_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na164_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na367_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a369_4 ( .OUT(na369_2), .COUTY1(na369_4), .IN1(1'b0), .IN2(1'b0), .IN3(na167_1), .IN4(1'b1), .IN5(na164_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na367_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y55     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a371_1 ( .OUT(na371_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na170_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na369_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a371_4 ( .OUT(na371_2), .COUTY1(na371_4), .IN1(1'b1), .IN2(na173_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na170_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na369_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y56     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a373_1 ( .OUT(na373_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na176_1),
                     .CINX(1'b0), .CINY1(na371_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a373_4 ( .OUT(na373_2), .COUTY1(na373_4), .IN1(na179_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na176_1), .CINX(1'b0), .CINY1(na371_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y57     80'h00_0078_00_0020_0C66_0AAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a375_1 ( .OUT(na375_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na182_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na373_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a375_4 ( .OUT(na375_2), .COUTY1(na375_4), .IN1(1'b1), .IN2(1'b1), .IN3(na186_1), .IN4(1'b1), .IN5(na182_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na373_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y58     80'h00_0078_00_0020_0C66_FAFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a378_1 ( .OUT(na378_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na189_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na375_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a378_4 ( .OUT(na378_2), .COUTY1(na378_4), .IN1(1'b1), .IN2(na193_1), .IN3(1'b1), .IN4(1'b1), .IN5(na189_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na375_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y59     80'h00_0078_00_0020_0C66_C0FA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a380_1 ( .OUT(na380_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na196_1),
                     .CINX(1'b0), .CINY1(na378_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a380_4 ( .OUT(na380_2), .COUTY1(na380_4), .IN1(na199_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na196_1), .CINX(1'b0), .CINY1(na378_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y60     80'h00_0078_00_0020_0C66_0AAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a382_1 ( .OUT(na382_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na202_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na380_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a382_4 ( .OUT(na382_2), .COUTY1(na382_4), .IN1(1'b1), .IN2(1'b1), .IN3(na205_1), .IN4(1'b1), .IN5(na202_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na380_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y61     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a384_1 ( .OUT(na384_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na315_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na382_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a384_4 ( .OUT(na384_2), .COUTY1(na384_4), .IN1(1'b1), .IN2(na209_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na315_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na382_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y62     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a386_1 ( .OUT(na386_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na212_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na384_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a386_4 ( .OUT(na386_2), .COUTY1(na386_4), .IN1(1'b1), .IN2(na215_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na212_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na384_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y35     80'h00_0078_00_0020_0C66_A0FA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a387_1 ( .OUT(na387_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na36_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na365_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a387_4 ( .OUT(na387_2), .COUTY1(na387_4), .IN1(na41_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na36_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na365_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y63     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a389_1 ( .OUT(na389_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na218_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na386_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a389_4 ( .OUT(na389_2), .IN1(na221_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na218_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na386_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y36     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a392_1 ( .OUT(na392_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na46_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na387_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a392_4 ( .OUT(na392_2), .COUTY1(na392_4), .IN1(1'b0), .IN2(1'b0), .IN3(na50_1), .IN4(1'b1), .IN5(1'b1), .IN6(na46_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na387_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x84y37     80'h00_0078_00_0020_0C66_CF0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a394_1 ( .OUT(na394_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na54_1),
                     .CINX(1'b0), .CINY1(na392_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a394_4 ( .OUT(na394_2), .COUTY1(na394_4), .IN1(1'b1), .IN2(na59_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na54_1), .CINX(1'b0), .CINY1(na392_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x84y32     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a395_2 ( .OUT(na395_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a395_6 ( .COUTY1(na395_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na395_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x86y40     80'h00_0078_00_0020_0C66_FCA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a397_1 ( .OUT(na397_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na59_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na458_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a397_4 ( .OUT(na397_2), .COUTY1(na397_4), .IN1(1'b0), .IN2(1'b0), .IN3(na62_1), .IN4(1'b1), .IN5(1'b1), .IN6(na59_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na458_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y41     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a399_1 ( .OUT(na399_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na66_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na397_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a399_4 ( .OUT(na399_2), .COUTY1(na399_4), .IN1(1'b0), .IN2(1'b0), .IN3(na69_1), .IN4(1'b1), .IN5(na66_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na397_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y42     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a401_1 ( .OUT(na401_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na72_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na399_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a401_4 ( .OUT(na401_2), .COUTY1(na401_4), .IN1(1'b0), .IN2(1'b0), .IN3(na75_1), .IN4(1'b1), .IN5(na72_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na399_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y43     80'h00_0078_00_0020_0C66_FCAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a403_1 ( .OUT(na403_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na78_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na401_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a403_4 ( .OUT(na403_2), .COUTY1(na403_4), .IN1(1'b1), .IN2(1'b1), .IN3(na81_1), .IN4(1'b1), .IN5(1'b1), .IN6(na78_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na401_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y44     80'h00_0078_00_0020_0C66_C0CF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a405_1 ( .OUT(na405_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na84_1),
                     .CINX(1'b0), .CINY1(na403_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a405_4 ( .OUT(na405_2), .COUTY1(na405_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na84_1), .CINX(1'b0), .CINY1(na403_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y35     80'h00_0078_00_0020_0C66_AACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a406_1 ( .OUT(na406_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na12_1), .IN6(1'b1), .IN7(na1_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na459_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a406_4 ( .OUT(na406_2), .COUTY1(na406_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na23_1), .IN5(na12_1), .IN6(1'b1), .IN7(na1_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na459_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y45     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a408_1 ( .OUT(na408_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na90_1),
                     .CINX(1'b0), .CINY1(na405_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a408_4 ( .OUT(na408_2), .COUTY1(na408_4), .IN1(na93_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na90_1), .CINX(1'b0), .CINY1(na405_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y46     80'h00_0078_00_0020_0C66_AF0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a410_1 ( .OUT(na410_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na96_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na408_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a410_4 ( .OUT(na410_2), .COUTY1(na410_4), .IN1(na99_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na96_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na408_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y47     80'h00_0078_00_0020_0C66_FAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a412_1 ( .OUT(na412_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na102_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na410_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a412_4 ( .OUT(na412_2), .COUTY1(na412_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na105_1), .IN5(na102_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na410_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y48     80'h00_0078_00_0020_0C66_0CAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a414_1 ( .OUT(na414_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na109_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na412_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a414_4 ( .OUT(na414_2), .COUTY1(na414_4), .IN1(1'b1), .IN2(1'b1), .IN3(na112_1), .IN4(1'b1), .IN5(1'b1), .IN6(na109_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na412_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y49     80'h00_0078_00_0020_0C66_FCAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a416_1 ( .OUT(na416_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na115_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na414_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a416_4 ( .OUT(na416_2), .COUTY1(na416_4), .IN1(1'b1), .IN2(1'b1), .IN3(na119_1), .IN4(1'b1), .IN5(1'b1), .IN6(na115_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na414_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y50     80'h00_0078_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a419_1 ( .OUT(na419_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na122_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na416_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a419_4 ( .OUT(na419_2), .COUTY1(na419_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na125_1), .IN5(1'b1), .IN6(na122_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na416_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y51     80'h00_0078_00_0020_0C66_FAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a421_1 ( .OUT(na421_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na128_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na419_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a421_4 ( .OUT(na421_2), .COUTY1(na421_4), .IN1(1'b0), .IN2(1'b0), .IN3(na131_1), .IN4(1'b1), .IN5(na128_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na419_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y52     80'h00_0078_00_0020_0C66_0AAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a423_1 ( .OUT(na423_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na134_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na421_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a423_4 ( .OUT(na423_2), .COUTY1(na423_4), .IN1(1'b1), .IN2(1'b1), .IN3(na137_1), .IN4(1'b1), .IN5(na134_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na421_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y53     80'h00_0078_00_0020_0C66_FCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a425_1 ( .OUT(na425_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na141_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na423_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a425_4 ( .OUT(na425_2), .COUTY1(na425_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na146_1), .IN5(1'b1), .IN6(na141_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na423_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y54     80'h00_0078_00_0020_0C66_FAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a427_1 ( .OUT(na427_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na149_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na425_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a427_4 ( .OUT(na427_2), .COUTY1(na427_4), .IN1(1'b1), .IN2(1'b1), .IN3(na152_1), .IN4(1'b1), .IN5(na149_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na425_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y36     80'h00_0078_00_0020_0C66_0AAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a428_1 ( .OUT(na428_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na27_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na406_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a428_4 ( .OUT(na428_2), .COUTY1(na428_4), .IN1(1'b1), .IN2(1'b1), .IN3(na30_1), .IN4(1'b1), .IN5(na27_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na406_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y55     80'h00_0078_00_0020_0C66_FCCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a430_1 ( .OUT(na430_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na155_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na427_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a430_4 ( .OUT(na430_2), .COUTY1(na430_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na158_1), .IN5(1'b1), .IN6(na155_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na427_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y56     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a432_1 ( .OUT(na432_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na161_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na430_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a432_4 ( .OUT(na432_2), .COUTY1(na432_4), .IN1(na164_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na161_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na430_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y57     80'h00_0078_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a434_1 ( .OUT(na434_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na167_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na432_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a434_4 ( .OUT(na434_2), .COUTY1(na434_4), .IN1(1'b1), .IN2(na170_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na167_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na432_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y58     80'h00_0078_00_0020_0C66_FCCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a436_1 ( .OUT(na436_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na173_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na434_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a436_4 ( .OUT(na436_2), .COUTY1(na436_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na176_1), .IN5(1'b1), .IN6(na173_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na434_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y59     80'h00_0078_00_0020_0C66_0AFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a438_1 ( .OUT(na438_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na179_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na436_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a438_4 ( .OUT(na438_2), .COUTY1(na438_4), .IN1(na182_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na179_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na436_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y60     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a441_1 ( .OUT(na441_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na186_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na438_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a441_4 ( .OUT(na441_2), .COUTY1(na441_4), .IN1(na189_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na186_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na438_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y61     80'h00_0078_00_0020_0C66_0CCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a443_1 ( .OUT(na443_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na193_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na441_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a443_4 ( .OUT(na443_2), .COUTY1(na443_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na196_1), .IN5(1'b1), .IN6(na193_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na441_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y62     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a445_1 ( .OUT(na445_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na199_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na443_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a445_4 ( .OUT(na445_2), .COUTY1(na445_4), .IN1(na202_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na199_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na443_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y63     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a447_1 ( .OUT(na447_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na205_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na445_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a447_4 ( .OUT(na447_2), .COUTY1(na447_4), .IN1(1'b0), .IN2(1'b0), .IN3(na315_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na205_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na445_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y64     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a449_1 ( .OUT(na449_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na209_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na447_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a449_4 ( .OUT(na449_2), .COUTY1(na449_4), .IN1(1'b0), .IN2(1'b0), .IN3(na212_1), .IN4(1'b1), .IN5(1'b1), .IN6(na209_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na447_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y37     80'h00_0078_00_0020_0C66_FAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a450_1 ( .OUT(na450_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na33_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na428_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a450_4 ( .OUT(na450_2), .COUTY1(na450_4), .IN1(1'b1), .IN2(1'b1), .IN3(na36_1), .IN4(1'b1), .IN5(na33_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na428_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y65     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a452_1 ( .OUT(na452_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na215_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na449_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a452_4 ( .OUT(na452_2), .COUTY1(na452_4), .IN1(1'b0), .IN2(1'b0), .IN3(na218_1), .IN4(1'b1), .IN5(1'b1), .IN6(na215_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na449_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x86y66     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a454_1 ( .OUT(na454_1), .IN1(na221_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na452_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y38     80'h00_0078_00_0020_0C66_0A0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a456_1 ( .OUT(na456_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na41_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na450_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a456_4 ( .OUT(na456_2), .COUTY1(na456_4), .IN1(1'b1), .IN2(na46_1), .IN3(1'b0), .IN4(1'b0), .IN5(na41_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na450_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x86y39     80'h00_0078_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a458_1 ( .OUT(na458_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na50_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na456_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a458_4 ( .OUT(na458_2), .COUTY1(na458_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na54_1), .IN5(1'b0), .IN6(1'b0), .IN7(na50_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na456_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x86y34     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a459_2 ( .OUT(na459_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a459_6 ( .COUTY1(na459_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na459_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x80y30     80'h00_EE60_00_0020_0C66_CCA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a460_1 ( .OUT(na460_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na789_1), .IN7(1'b1), .IN8(na460_1),
                     .CINX(1'b0), .CINY1(na462_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a460_2 ( .OUT(na460_1), .CLK(na685_1), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na460_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a460_4 ( .OUT(na460_2), .IN1(1'b0), .IN2(1'b0), .IN3(na685_3), .IN4(1'b1), .IN5(1'b1), .IN6(na789_1), .IN7(1'b1), .IN8(na460_1),
                     .CINX(1'b0), .CINY1(na462_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x80y29     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a462_2 ( .OUT(na462_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a462_6 ( .COUTY1(na462_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na462_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x79y59     80'h00_ED60_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a463_1 ( .OUT(na463_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na463_1), .IN6(1'b1), .IN7(1'b1), .IN8(na780_1),
                     .CINX(1'b0), .CINY1(na532_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a463_2 ( .OUT(na463_1), .CLK(~na685_3), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na463_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a463_4 ( .OUT(na463_2), .COUTY1(na463_4), .IN1(na782_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na463_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na780_1), .CINX(1'b0), .CINY1(na532_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x79y60     80'h00_ED60_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a465_1 ( .OUT(na465_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na465_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na463_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a465_2 ( .OUT(na465_1), .CLK(~na685_3), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na465_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a465_4 ( .OUT(na465_2), .COUTY1(na465_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na784_1), .IN5(1'b1), .IN6(na465_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na463_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF/D///      x79y61     80'h00_ED00_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a467_1 ( .OUT(na467_1_i), .IN1(1'b1), .IN2(na685_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na465_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a467_2 ( .OUT(na467_1), .CLK(~na685_3), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na467_1_i) );
// C_ADDF2/D//ADDF2/      x87y34     80'h00_EE60_00_0020_0C66_ACAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a468_1 ( .OUT(na468_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na468_1), .IN7(na1_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na535_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a468_2 ( .OUT(na468_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na468_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a468_4 ( .OUT(na468_2), .COUTY1(na468_4), .IN1(na12_1), .IN2(1'b1), .IN3(na717_2), .IN4(1'b1), .IN5(1'b1), .IN6(na468_1),
                     .IN7(na1_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na535_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y39     80'h00_EE60_00_0020_0C66_CACC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a469_1 ( .OUT(na469_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na469_1), .IN6(1'b1), .IN7(1'b1), .IN8(na54_1),
                     .CINX(1'b0), .CINY1(na530_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a469_2 ( .OUT(na469_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na469_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a469_4 ( .OUT(na469_2), .COUTY1(na469_4), .IN1(1'b1), .IN2(na59_1), .IN3(1'b1), .IN4(na727_1), .IN5(na469_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na54_1), .CINX(1'b0), .CINY1(na530_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y40     80'h00_EE60_00_0020_0C66_ACAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a471_1 ( .OUT(na471_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na471_1), .IN7(na62_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na469_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a471_2 ( .OUT(na471_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na471_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a471_4 ( .OUT(na471_2), .COUTY1(na471_4), .IN1(na66_1), .IN2(1'b1), .IN3(na729_2), .IN4(1'b1), .IN5(1'b1), .IN6(na471_1),
                     .IN7(na62_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na469_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y41     80'h00_EE60_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a473_1 ( .OUT(na473_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na473_1), .IN6(1'b1), .IN7(na69_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na471_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a473_2 ( .OUT(na473_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na473_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a473_4 ( .OUT(na473_2), .COUTY1(na473_4), .IN1(na72_1), .IN2(1'b1), .IN3(na731_1), .IN4(1'b1), .IN5(na473_1), .IN6(1'b1),
                     .IN7(na69_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na471_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y42     80'h00_EE60_00_0020_0C66_ACAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a475_1 ( .OUT(na475_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na475_1), .IN7(na75_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na473_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a475_2 ( .OUT(na475_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na475_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a475_4 ( .OUT(na475_2), .COUTY1(na475_4), .IN1(1'b1), .IN2(na78_1), .IN3(na733_1), .IN4(1'b1), .IN5(1'b1), .IN6(na475_1),
                     .IN7(na75_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na473_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y43     80'h00_EE60_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a477_1 ( .OUT(na477_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na477_1), .IN6(1'b1), .IN7(na81_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na475_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a477_2 ( .OUT(na477_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na477_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a477_4 ( .OUT(na477_2), .COUTY1(na477_4), .IN1(na735_1), .IN2(1'b1), .IN3(1'b1), .IN4(na84_1), .IN5(na477_1), .IN6(1'b1),
                     .IN7(na81_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na475_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y44     80'h00_EE60_00_0020_0C66_CCCC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a480_1 ( .OUT(na480_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na480_1), .IN7(1'b1), .IN8(na87_1),
                     .CINX(1'b0), .CINY1(na477_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a480_2 ( .OUT(na480_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na480_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a480_4 ( .OUT(na480_2), .COUTY1(na480_4), .IN1(1'b1), .IN2(na737_2), .IN3(1'b1), .IN4(na90_1), .IN5(1'b1), .IN6(na480_1),
                     .IN7(1'b1), .IN8(na87_1), .CINX(1'b0), .CINY1(na477_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y45     80'h00_EE60_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a482_1 ( .OUT(na482_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na482_1), .IN6(1'b1), .IN7(na1234_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na480_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a482_2 ( .OUT(na482_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na482_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a482_4 ( .OUT(na482_2), .COUTY1(na482_4), .IN1(na739_1), .IN2(1'b1), .IN3(na96_1), .IN4(1'b1), .IN5(na482_1), .IN6(1'b1),
                     .IN7(na1234_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na480_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y46     80'h00_EE60_00_0020_0C66_ACAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a484_1 ( .OUT(na484_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na484_1), .IN7(na1235_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na482_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a484_2 ( .OUT(na484_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na484_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a484_4 ( .OUT(na484_2), .COUTY1(na484_4), .IN1(na102_1), .IN2(1'b1), .IN3(na741_2), .IN4(1'b1), .IN5(1'b1), .IN6(na484_1),
                     .IN7(na1235_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na482_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y47     80'h00_EE60_00_0020_0C66_CAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a486_1 ( .OUT(na486_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na486_1), .IN6(1'b1), .IN7(1'b1), .IN8(na105_1),
                     .CINX(1'b0), .CINY1(na484_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a486_2 ( .OUT(na486_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na486_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a486_4 ( .OUT(na486_2), .COUTY1(na486_4), .IN1(1'b1), .IN2(na109_1), .IN3(na743_2), .IN4(1'b1), .IN5(na486_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na105_1), .CINX(1'b0), .CINY1(na484_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y48     80'h00_EE60_00_0020_0C66_ACAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a488_1 ( .OUT(na488_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na488_1), .IN7(na112_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na486_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a488_2 ( .OUT(na488_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na488_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a488_4 ( .OUT(na488_2), .COUTY1(na488_4), .IN1(1'b1), .IN2(na115_1), .IN3(na745_2), .IN4(1'b1), .IN5(1'b1), .IN6(na488_1),
                     .IN7(na112_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na486_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y35     80'h00_EE60_00_0020_0C66_CAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a490_1 ( .OUT(na490_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na490_1), .IN6(1'b1), .IN7(1'b1), .IN8(na23_1),
                     .CINX(1'b0), .CINY1(na468_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a490_2 ( .OUT(na490_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na490_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a490_4 ( .OUT(na490_2), .COUTY1(na490_4), .IN1(na27_1), .IN2(1'b1), .IN3(na719_1), .IN4(1'b1), .IN5(na490_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na23_1), .CINX(1'b0), .CINY1(na468_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y49     80'h00_EE60_00_0020_0C66_AAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a491_1 ( .OUT(na491_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na491_1), .IN6(1'b1), .IN7(na119_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na488_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a491_2 ( .OUT(na491_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na491_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a491_4 ( .OUT(na491_2), .COUTY1(na491_4), .IN1(1'b1), .IN2(na122_1), .IN3(na747_1), .IN4(1'b1), .IN5(na491_1), .IN6(1'b1),
                     .IN7(na119_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na488_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y50     80'h00_EE60_00_0020_0C66_CCAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a493_1 ( .OUT(na493_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na493_1), .IN7(1'b1), .IN8(na125_1),
                     .CINX(1'b0), .CINY1(na491_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a493_2 ( .OUT(na493_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na493_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a493_4 ( .OUT(na493_2), .COUTY1(na493_4), .IN1(na128_1), .IN2(1'b1), .IN3(na749_1), .IN4(1'b1), .IN5(1'b1), .IN6(na493_1),
                     .IN7(1'b1), .IN8(na125_1), .CINX(1'b0), .CINY1(na491_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y51     80'h00_EE60_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a495_1 ( .OUT(na495_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na495_1), .IN6(1'b1), .IN7(na131_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na493_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a495_2 ( .OUT(na495_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na495_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a495_4 ( .OUT(na495_2), .COUTY1(na495_4), .IN1(na134_1), .IN2(1'b1), .IN3(1'b1), .IN4(na751_1), .IN5(na495_1), .IN6(1'b1),
                     .IN7(na131_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na493_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y52     80'h00_EE60_00_0020_0C66_ACAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a497_1 ( .OUT(na497_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na497_1), .IN7(na137_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na495_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a497_2 ( .OUT(na497_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na497_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a497_4 ( .OUT(na497_2), .COUTY1(na497_4), .IN1(1'b1), .IN2(na141_1), .IN3(na753_2), .IN4(1'b1), .IN5(1'b1), .IN6(na497_1),
                     .IN7(na137_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na495_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y53     80'h00_EE60_00_0020_0C66_CAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a499_1 ( .OUT(na499_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na499_1), .IN6(1'b1), .IN7(1'b1), .IN8(na146_1),
                     .CINX(1'b0), .CINY1(na497_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a499_2 ( .OUT(na499_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na499_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a499_4 ( .OUT(na499_2), .COUTY1(na499_4), .IN1(na149_1), .IN2(1'b1), .IN3(na755_2), .IN4(1'b1), .IN5(na499_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na146_1), .CINX(1'b0), .CINY1(na497_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y54     80'h00_EE60_00_0020_0C66_ACAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a502_1 ( .OUT(na502_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na502_1), .IN7(na152_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na499_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a502_2 ( .OUT(na502_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na502_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a502_4 ( .OUT(na502_2), .COUTY1(na502_4), .IN1(1'b1), .IN2(na155_1), .IN3(na757_2), .IN4(1'b1), .IN5(1'b1), .IN6(na502_1),
                     .IN7(na152_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na499_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y55     80'h00_EE60_00_0020_0C66_CACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a504_1 ( .OUT(na504_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na504_1), .IN6(1'b1), .IN7(1'b1), .IN8(na158_1),
                     .CINX(1'b0), .CINY1(na502_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a504_2 ( .OUT(na504_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na504_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a504_4 ( .OUT(na504_2), .COUTY1(na504_4), .IN1(na161_1), .IN2(1'b1), .IN3(1'b1), .IN4(na759_1), .IN5(na504_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na158_1), .CINX(1'b0), .CINY1(na502_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y56     80'h00_EE60_00_0020_0C66_ACAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a506_1 ( .OUT(na506_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na506_1), .IN7(na1237_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na504_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a506_2 ( .OUT(na506_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na506_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a506_4 ( .OUT(na506_2), .COUTY1(na506_4), .IN1(1'b1), .IN2(na761_2), .IN3(na167_1), .IN4(1'b1), .IN5(1'b1), .IN6(na506_1),
                     .IN7(na1237_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na504_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y57     80'h00_EE60_00_0020_0C66_CACC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a508_1 ( .OUT(na508_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na508_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1238_2),
                     .CINX(1'b0), .CINY1(na506_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a508_2 ( .OUT(na508_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na508_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a508_4 ( .OUT(na508_2), .COUTY1(na508_4), .IN1(1'b1), .IN2(na173_1), .IN3(1'b1), .IN4(na763_1), .IN5(na508_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na1238_2), .CINX(1'b0), .CINY1(na506_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y58     80'h00_EE60_00_0020_0C66_CCAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a510_1 ( .OUT(na510_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na510_1), .IN7(1'b1), .IN8(na176_1),
                     .CINX(1'b0), .CINY1(na508_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a510_2 ( .OUT(na510_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na510_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a510_4 ( .OUT(na510_2), .COUTY1(na510_4), .IN1(na179_1), .IN2(1'b1), .IN3(na765_1), .IN4(1'b1), .IN5(1'b1), .IN6(na510_1),
                     .IN7(1'b1), .IN8(na176_1), .CINX(1'b0), .CINY1(na508_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y36     80'h00_EE60_00_0020_0C66_ACAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a512_1 ( .OUT(na512_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na512_1), .IN7(na30_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na490_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a512_2 ( .OUT(na512_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na512_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a512_4 ( .OUT(na512_2), .COUTY1(na512_4), .IN1(na33_1), .IN2(1'b1), .IN3(na721_2), .IN4(1'b1), .IN5(1'b1), .IN6(na512_1),
                     .IN7(na30_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na490_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y59     80'h00_EE60_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a513_1 ( .OUT(na513_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na513_1), .IN6(1'b1), .IN7(na1239_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na510_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a513_2 ( .OUT(na513_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na513_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a513_4 ( .OUT(na513_2), .COUTY1(na513_4), .IN1(na767_1), .IN2(1'b1), .IN3(na186_1), .IN4(1'b1), .IN5(na513_1), .IN6(1'b1),
                     .IN7(na1239_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na510_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y60     80'h00_EE60_00_0020_0C66_ACCC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a515_1 ( .OUT(na515_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na515_1), .IN7(na1240_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na513_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a515_2 ( .OUT(na515_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na515_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a515_4 ( .OUT(na515_2), .COUTY1(na515_4), .IN1(1'b1), .IN2(na193_1), .IN3(1'b1), .IN4(na769_2), .IN5(1'b1), .IN6(na515_1),
                     .IN7(na1240_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na513_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y61     80'h00_EE60_00_0020_0C66_CAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a517_1 ( .OUT(na517_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na517_1), .IN6(1'b1), .IN7(1'b1), .IN8(na196_1),
                     .CINX(1'b0), .CINY1(na515_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a517_2 ( .OUT(na517_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na517_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a517_4 ( .OUT(na517_2), .COUTY1(na517_4), .IN1(na199_1), .IN2(1'b1), .IN3(na771_1), .IN4(1'b1), .IN5(na517_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na196_1), .CINX(1'b0), .CINY1(na515_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y62     80'h00_EE60_00_0020_0C66_ACAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a519_1 ( .OUT(na519_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na519_1), .IN7(na1241_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na517_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a519_2 ( .OUT(na519_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na519_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a519_4 ( .OUT(na519_2), .COUTY1(na519_4), .IN1(1'b1), .IN2(na773_2), .IN3(na205_1), .IN4(1'b1), .IN5(1'b1), .IN6(na519_1),
                     .IN7(na1241_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na517_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y63     80'h00_EE60_00_0020_0C66_AAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a521_1 ( .OUT(na521_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na521_1), .IN6(1'b1), .IN7(na315_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na519_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a521_2 ( .OUT(na521_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na521_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a521_4 ( .OUT(na521_2), .COUTY1(na521_4), .IN1(1'b1), .IN2(na209_1), .IN3(na775_2), .IN4(1'b1), .IN5(na521_1), .IN6(1'b1),
                     .IN7(na315_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na519_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y64     80'h00_EE60_00_0020_0C66_ACAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a524_1 ( .OUT(na524_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na524_1), .IN7(na212_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na521_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a524_2 ( .OUT(na524_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na524_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a524_4 ( .OUT(na524_2), .COUTY1(na524_4), .IN1(1'b1), .IN2(na215_1), .IN3(na777_2), .IN4(1'b1), .IN5(1'b1), .IN6(na524_1),
                     .IN7(na212_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na521_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y65     80'h00_EE60_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a526_1 ( .OUT(na526_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na526_1), .IN6(1'b1), .IN7(na218_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na524_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a526_2 ( .OUT(na526_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na526_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a526_4 ( .OUT(na526_2), .IN1(na221_1), .IN2(1'b1), .IN3(na779_1), .IN4(1'b1), .IN5(na526_1), .IN6(1'b1), .IN7(na218_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na524_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y37     80'h00_EE60_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a528_1 ( .OUT(na528_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na528_1), .IN6(1'b1), .IN7(na36_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na512_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a528_2 ( .OUT(na528_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na528_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a528_4 ( .OUT(na528_2), .COUTY1(na528_4), .IN1(na41_1), .IN2(1'b1), .IN3(1'b1), .IN4(na723_2), .IN5(na528_1), .IN6(1'b1),
                     .IN7(na36_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na512_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x87y38     80'h00_EE60_00_0020_0C66_CCAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a530_1 ( .OUT(na530_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na530_1), .IN7(1'b1), .IN8(na1232_2),
                     .CINX(1'b0), .CINY1(na528_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a530_2 ( .OUT(na530_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na530_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a530_4 ( .OUT(na530_2), .COUTY1(na530_4), .IN1(na725_2), .IN2(1'b1), .IN3(na50_1), .IN4(1'b1), .IN5(1'b1), .IN6(na530_1),
                     .IN7(1'b1), .IN8(na1232_2), .CINX(1'b0), .CINY1(na528_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x79y58     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a532_2 ( .OUT(na532_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a532_6 ( .COUTY1(na532_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na532_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x82y31     80'h00_0078_00_0020_0C66_AA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a533_1 ( .OUT(na533_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na265_2), .IN6(1'b1), .IN7(na1249_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na551_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a533_4 ( .OUT(na533_2), .IN1(1'b1), .IN2(na262_1), .IN3(1'b0), .IN4(1'b0), .IN5(na265_2), .IN6(1'b1), .IN7(na1249_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na551_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x87y33     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a535_2 ( .OUT(na535_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a535_6 ( .COUTY1(na535_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na535_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x92y36     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a537_1 ( .OUT(na537_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na246_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na550_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a537_4 ( .OUT(na537_2), .COUTY1(na537_4), .IN1(na247_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na246_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na550_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x92y37     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a539_1 ( .OUT(na539_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na247_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na537_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a539_4 ( .OUT(na539_2), .COUTY1(na539_4), .IN1(1'b0), .IN2(1'b0), .IN3(na249_2), .IN4(1'b1), .IN5(na247_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na537_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x92y38     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a541_1 ( .OUT(na541_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na250_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na539_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x92y31     80'h00_0078_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a542_1 ( .OUT(na542_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na236_1), .IN7(1'b1), .IN8(na237_2),
                     .CINX(1'b0), .CINY1(na554_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a542_4 ( .OUT(na542_2), .COUTY1(na542_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na237_1), .IN5(1'b1), .IN6(na236_1), .IN7(1'b1),
                     .IN8(na237_2), .CINX(1'b0), .CINY1(na554_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x92y32     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a544_1 ( .OUT(na544_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na239_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na542_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a544_4 ( .OUT(na544_2), .COUTY1(na544_4), .IN1(na239_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na239_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na542_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x92y33     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a546_1 ( .OUT(na546_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na241_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na544_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a546_4 ( .OUT(na546_2), .COUTY1(na546_4), .IN1(1'b1), .IN2(na241_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na241_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na544_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x92y34     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a548_1 ( .OUT(na548_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na243_2),
                     .CINX(1'b0), .CINY1(na546_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a548_4 ( .OUT(na548_2), .COUTY1(na548_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na243_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na243_2), .CINX(1'b0), .CINY1(na546_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x92y35     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a550_1 ( .OUT(na550_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na245_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na548_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a550_4 ( .OUT(na550_2), .COUTY1(na550_4), .IN1(1'b1), .IN2(na245_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na245_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na548_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x82y30     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a551_2 ( .OUT(na551_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a551_6 ( .COUTY1(na551_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na551_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x84y30     80'h00_0078_00_0020_0C66_5503
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a552_1 ( .OUT(na552_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na265_2), .IN6(1'b1), .IN7(~na1249_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na555_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a552_4 ( .OUT(na552_2), .COUTY1(na552_4), .IN1(1'b1), .IN2(~na262_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na265_2), .IN6(1'b1),
                     .IN7(~na1249_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na555_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x92y30     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a554_2 ( .OUT(na554_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a554_6 ( .COUTY1(na554_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na554_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x84y29     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a555_2 ( .OUT(na555_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a555_6 ( .COUTY1(na555_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na555_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x88y40     80'h00_0078_00_0020_0C66_A0FA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a557_1 ( .OUT(na557_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(na62_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na617_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a557_4 ( .OUT(na557_2), .COUTY1(na557_4), .IN1(na66_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(na62_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na617_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y41     80'h00_0078_00_0020_0C66_A0FA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a559_1 ( .OUT(na559_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(na69_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na557_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a559_4 ( .OUT(na559_2), .COUTY1(na559_4), .IN1(na72_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(na69_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na557_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y42     80'h00_0078_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a561_1 ( .OUT(na561_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na75_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na559_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a561_4 ( .OUT(na561_2), .COUTY1(na561_4), .IN1(1'b1), .IN2(na78_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na75_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na559_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y43     80'h00_0078_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a563_1 ( .OUT(na563_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(na81_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na561_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a563_4 ( .OUT(na563_2), .COUTY1(na563_4), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(na84_1), .IN5(1'b0), .IN6(1'b1), .IN7(na81_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na561_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y44     80'h00_0078_00_0020_0C66_C0CF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a565_1 ( .OUT(na565_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(na87_1),
                     .CINX(1'b0), .CINY1(na563_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a565_4 ( .OUT(na565_2), .COUTY1(na565_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na90_1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na87_1), .CINX(1'b0), .CINY1(na563_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y35     80'h00_0078_00_0020_0C66_CAFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a566_1 ( .OUT(na566_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na12_1), .IN6(1'b1), .IN7(1'b1), .IN8(na23_1),
                     .CINX(1'b0), .CINY1(na618_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a566_4 ( .OUT(na566_2), .COUTY1(na566_4), .IN1(na27_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na12_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na23_1), .CINX(1'b0), .CINY1(na618_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y45     80'h00_0078_00_0020_0C66_FAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a568_1 ( .OUT(na568_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na93_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na565_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a568_4 ( .OUT(na568_2), .COUTY1(na568_4), .IN1(1'b0), .IN2(1'b1), .IN3(na96_1), .IN4(1'b1), .IN5(na93_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na565_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y46     80'h00_0078_00_0020_0C66_0AFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a570_1 ( .OUT(na570_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na99_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na568_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a570_4 ( .OUT(na570_2), .COUTY1(na570_4), .IN1(na102_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na99_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na568_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y47     80'h00_0078_00_0020_0C66_C00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a572_1 ( .OUT(na572_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(na105_1),
                     .CINX(1'b0), .CINY1(na570_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a572_4 ( .OUT(na572_2), .COUTY1(na572_4), .IN1(1'b1), .IN2(na109_1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na105_1), .CINX(1'b0), .CINY1(na570_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y48     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a574_1 ( .OUT(na574_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(na112_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na572_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a574_4 ( .OUT(na574_2), .COUTY1(na574_4), .IN1(1'b1), .IN2(na115_1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(na112_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na572_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y49     80'h00_0078_00_0020_0C66_A0FC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a576_1 ( .OUT(na576_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(na119_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na574_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a576_4 ( .OUT(na576_2), .COUTY1(na576_4), .IN1(1'b1), .IN2(na122_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(na119_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na574_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y50     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a579_1 ( .OUT(na579_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na125_1),
                     .CINX(1'b0), .CINY1(na576_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a579_4 ( .OUT(na579_2), .COUTY1(na579_4), .IN1(na128_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na125_1), .CINX(1'b0), .CINY1(na576_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y51     80'h00_0078_00_0020_0C66_AF0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a581_1 ( .OUT(na581_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na131_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na579_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a581_4 ( .OUT(na581_2), .COUTY1(na581_4), .IN1(na134_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na131_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na579_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y52     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a583_1 ( .OUT(na583_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(na137_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na581_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a583_4 ( .OUT(na583_2), .COUTY1(na583_4), .IN1(1'b1), .IN2(na141_1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(na137_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na581_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y53     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a585_1 ( .OUT(na585_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(na146_1),
                     .CINX(1'b0), .CINY1(na583_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a585_4 ( .OUT(na585_2), .COUTY1(na585_4), .IN1(na149_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na146_1), .CINX(1'b0), .CINY1(na583_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y54     80'h00_0078_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a587_1 ( .OUT(na587_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na152_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na585_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a587_4 ( .OUT(na587_2), .COUTY1(na587_4), .IN1(1'b1), .IN2(na155_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na152_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na585_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y36     80'h00_0078_00_0020_0C66_AF0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a588_1 ( .OUT(na588_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na30_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na566_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a588_4 ( .OUT(na588_2), .COUTY1(na588_4), .IN1(na33_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na30_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na566_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y55     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a590_1 ( .OUT(na590_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(na158_1),
                     .CINX(1'b0), .CINY1(na587_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a590_4 ( .OUT(na590_2), .COUTY1(na590_4), .IN1(na161_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na158_1), .CINX(1'b0), .CINY1(na587_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y56     80'h00_0078_00_0020_0C66_FAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a592_1 ( .OUT(na592_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na164_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na590_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a592_4 ( .OUT(na592_2), .COUTY1(na592_4), .IN1(1'b1), .IN2(1'b1), .IN3(na167_1), .IN4(1'b1), .IN5(na164_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na590_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y57     80'h00_0078_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a594_1 ( .OUT(na594_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na170_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na592_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a594_4 ( .OUT(na594_2), .COUTY1(na594_4), .IN1(1'b1), .IN2(na173_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na170_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na592_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y58     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a596_1 ( .OUT(na596_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(na176_1),
                     .CINX(1'b0), .CINY1(na594_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a596_4 ( .OUT(na596_2), .COUTY1(na596_4), .IN1(na179_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na176_1), .CINX(1'b0), .CINY1(na594_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y59     80'h00_0078_00_0020_0C66_FAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a598_1 ( .OUT(na598_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na182_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na596_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a598_4 ( .OUT(na598_2), .COUTY1(na598_4), .IN1(1'b0), .IN2(1'b1), .IN3(na186_1), .IN4(1'b1), .IN5(na182_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na596_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y60     80'h00_0078_00_0020_0C66_0A0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a601_1 ( .OUT(na601_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na189_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na598_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a601_4 ( .OUT(na601_2), .COUTY1(na601_4), .IN1(1'b1), .IN2(na193_1), .IN3(1'b0), .IN4(1'b1), .IN5(na189_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na598_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y61     80'h00_0078_00_0020_0C66_CF0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a603_1 ( .OUT(na603_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na196_1),
                     .CINX(1'b0), .CINY1(na601_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a603_4 ( .OUT(na603_2), .COUTY1(na603_4), .IN1(na199_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na196_1), .CINX(1'b0), .CINY1(na601_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y62     80'h00_0078_00_0020_0C66_FAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a605_1 ( .OUT(na605_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na202_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na603_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a605_4 ( .OUT(na605_2), .COUTY1(na605_4), .IN1(1'b0), .IN2(1'b1), .IN3(na205_1), .IN4(1'b1), .IN5(na202_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na603_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y63     80'h00_0078_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a607_1 ( .OUT(na607_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na315_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na605_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a607_4 ( .OUT(na607_2), .COUTY1(na607_4), .IN1(1'b1), .IN2(na209_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na315_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na605_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y64     80'h00_0078_00_0020_0C66_AFFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a609_1 ( .OUT(na609_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na212_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na607_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a609_4 ( .OUT(na609_2), .COUTY1(na609_4), .IN1(1'b1), .IN2(na215_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na212_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na607_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y37     80'h00_0078_00_0020_0C66_AF0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a610_1 ( .OUT(na610_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na36_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na588_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a610_4 ( .OUT(na610_2), .COUTY1(na610_4), .IN1(na41_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na36_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na588_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y65     80'h00_0078_00_0020_0C66_AFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a612_1 ( .OUT(na612_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na218_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na609_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a612_4 ( .OUT(na612_2), .IN1(na221_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na218_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na609_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y38     80'h00_0078_00_0020_0C66_FCAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a615_1 ( .OUT(na615_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na46_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na610_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a615_4 ( .OUT(na615_2), .COUTY1(na615_4), .IN1(1'b1), .IN2(1'b1), .IN3(na50_1), .IN4(1'b1), .IN5(1'b1), .IN6(na46_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na610_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x88y39     80'h00_0078_00_0020_0C66_C0FC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a617_1 ( .OUT(na617_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(na54_1),
                     .CINX(1'b0), .CINY1(na615_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a617_4 ( .OUT(na617_2), .COUTY1(na617_4), .IN1(1'b1), .IN2(na59_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na54_1), .CINX(1'b0), .CINY1(na615_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x88y34     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a618_2 ( .OUT(na618_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a618_6 ( .COUTY1(na618_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na618_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x85y40     80'h00_0078_00_0020_0C66_0CAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a620_1 ( .OUT(na620_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na59_1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na681_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a620_4 ( .OUT(na620_2), .COUTY1(na620_4), .IN1(1'b1), .IN2(1'b1), .IN3(na62_1), .IN4(1'b1), .IN5(1'b1), .IN6(na59_1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na681_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y41     80'h00_0078_00_0020_0C66_FAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a622_1 ( .OUT(na622_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na66_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na620_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a622_4 ( .OUT(na622_2), .COUTY1(na622_4), .IN1(1'b1), .IN2(1'b1), .IN3(na69_1), .IN4(1'b1), .IN5(na66_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na620_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y42     80'h00_0078_00_0020_0C66_FAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a624_1 ( .OUT(na624_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na72_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na622_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a624_4 ( .OUT(na624_2), .COUTY1(na624_4), .IN1(1'b1), .IN2(1'b1), .IN3(na75_1), .IN4(1'b1), .IN5(na72_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na622_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y43     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a626_1 ( .OUT(na626_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na78_1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na624_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a626_4 ( .OUT(na626_2), .COUTY1(na626_4), .IN1(1'b0), .IN2(1'b1), .IN3(na81_1), .IN4(1'b1), .IN5(1'b1), .IN6(na78_1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na624_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y44     80'h00_0078_00_0020_0C66_CFC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a628_1 ( .OUT(na628_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na84_1),
                     .CINX(1'b0), .CINY1(na626_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a628_4 ( .OUT(na628_2), .COUTY1(na628_4), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na84_1), .CINX(1'b0), .CINY1(na626_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y35     80'h00_0078_00_0020_0C66_AAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a629_1 ( .OUT(na629_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na12_1), .IN6(1'b1), .IN7(na1_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na898_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a629_4 ( .OUT(na629_2), .COUTY1(na629_4), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(na23_1), .IN5(na12_1), .IN6(1'b1), .IN7(na1_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na898_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y45     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a631_1 ( .OUT(na631_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(na90_1),
                     .CINX(1'b0), .CINY1(na628_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a631_4 ( .OUT(na631_2), .COUTY1(na631_4), .IN1(na93_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na90_1), .CINX(1'b0), .CINY1(na628_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y46     80'h00_0078_00_0020_0C66_A0FA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a633_1 ( .OUT(na633_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(na96_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na631_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a633_4 ( .OUT(na633_2), .COUTY1(na633_4), .IN1(na99_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(na96_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na631_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y47     80'h00_0078_00_0020_0C66_0ACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a635_1 ( .OUT(na635_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na102_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na633_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a635_4 ( .OUT(na635_2), .COUTY1(na635_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na105_1), .IN5(na102_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na633_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y48     80'h00_0078_00_0020_0C66_FCA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a637_1 ( .OUT(na637_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na109_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na635_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a637_4 ( .OUT(na637_2), .COUTY1(na637_4), .IN1(1'b0), .IN2(1'b1), .IN3(na112_1), .IN4(1'b1), .IN5(1'b1), .IN6(na109_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na635_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y49     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a639_1 ( .OUT(na639_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na115_1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na637_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a639_4 ( .OUT(na639_2), .COUTY1(na639_4), .IN1(1'b0), .IN2(1'b1), .IN3(na119_1), .IN4(1'b1), .IN5(1'b1), .IN6(na115_1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na637_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y50     80'h00_0078_00_0020_0C66_FCCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a642_1 ( .OUT(na642_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na122_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na639_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a642_4 ( .OUT(na642_2), .COUTY1(na642_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na125_1), .IN5(1'b1), .IN6(na122_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na639_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y51     80'h00_0078_00_0020_0C66_0AAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a644_1 ( .OUT(na644_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na128_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na642_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a644_4 ( .OUT(na644_2), .COUTY1(na644_4), .IN1(1'b1), .IN2(1'b1), .IN3(na131_1), .IN4(1'b1), .IN5(na128_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na642_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y52     80'h00_0078_00_0020_0C66_FAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a646_1 ( .OUT(na646_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na134_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na644_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a646_4 ( .OUT(na646_2), .COUTY1(na646_4), .IN1(1'b0), .IN2(1'b1), .IN3(na137_1), .IN4(1'b1), .IN5(na134_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na644_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y53     80'h00_0078_00_0020_0C66_0CCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a648_1 ( .OUT(na648_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na141_1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na646_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a648_4 ( .OUT(na648_2), .COUTY1(na648_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na146_1), .IN5(1'b1), .IN6(na141_1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na646_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y54     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a650_1 ( .OUT(na650_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na149_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na648_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a650_4 ( .OUT(na650_2), .COUTY1(na650_4), .IN1(1'b0), .IN2(1'b1), .IN3(na152_1), .IN4(1'b1), .IN5(na149_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na648_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y36     80'h00_0078_00_0020_0C66_FAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a651_1 ( .OUT(na651_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na27_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na629_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a651_4 ( .OUT(na651_2), .COUTY1(na651_4), .IN1(1'b0), .IN2(1'b1), .IN3(na30_1), .IN4(1'b1), .IN5(na27_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na629_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y55     80'h00_0078_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a653_1 ( .OUT(na653_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na155_1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na650_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a653_4 ( .OUT(na653_2), .COUTY1(na653_4), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(na158_1), .IN5(1'b1), .IN6(na155_1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na650_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y56     80'h00_0078_00_0020_0C66_FAFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a655_1 ( .OUT(na655_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na161_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na653_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a655_4 ( .OUT(na655_2), .COUTY1(na655_4), .IN1(na164_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na161_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na653_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y57     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a657_1 ( .OUT(na657_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(na167_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na655_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a657_4 ( .OUT(na657_2), .COUTY1(na657_4), .IN1(1'b1), .IN2(na170_1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(na167_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na655_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y58     80'h00_0078_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a659_1 ( .OUT(na659_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na173_1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na657_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a659_4 ( .OUT(na659_2), .COUTY1(na659_4), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(na176_1), .IN5(1'b1), .IN6(na173_1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na657_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y59     80'h00_0078_00_0020_0C66_FA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a661_1 ( .OUT(na661_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na179_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na659_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a661_4 ( .OUT(na661_2), .COUTY1(na661_4), .IN1(na182_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b1), .IN5(na179_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na659_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y60     80'h00_0078_00_0020_0C66_AFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a664_1 ( .OUT(na664_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na186_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na661_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a664_4 ( .OUT(na664_2), .COUTY1(na664_4), .IN1(na189_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na186_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na661_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y61     80'h00_0078_00_0020_0C66_FCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a666_1 ( .OUT(na666_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na193_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na664_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a666_4 ( .OUT(na666_2), .COUTY1(na666_4), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(na196_1), .IN5(1'b1), .IN6(na193_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na664_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y62     80'h00_0078_00_0020_0C66_FAFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a668_1 ( .OUT(na668_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na199_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na666_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a668_4 ( .OUT(na668_2), .COUTY1(na668_4), .IN1(na202_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na199_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na666_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y63     80'h00_0078_00_0020_0C66_AFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a670_1 ( .OUT(na670_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na205_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na668_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a670_4 ( .OUT(na670_2), .COUTY1(na670_4), .IN1(1'b1), .IN2(1'b1), .IN3(na315_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na205_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na668_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y64     80'h00_0078_00_0020_0C66_FCAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a672_1 ( .OUT(na672_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na209_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na670_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a672_4 ( .OUT(na672_2), .COUTY1(na672_4), .IN1(1'b1), .IN2(1'b1), .IN3(na212_1), .IN4(1'b1), .IN5(1'b1), .IN6(na209_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na670_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y37     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a673_1 ( .OUT(na673_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na33_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na651_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a673_4 ( .OUT(na673_2), .COUTY1(na673_4), .IN1(1'b0), .IN2(1'b1), .IN3(na36_1), .IN4(1'b1), .IN5(na33_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na651_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y65     80'h00_0078_00_0020_0C66_FCAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a675_1 ( .OUT(na675_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na215_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na672_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a675_4 ( .OUT(na675_2), .COUTY1(na675_4), .IN1(1'b1), .IN2(1'b1), .IN3(na218_1), .IN4(1'b1), .IN5(1'b1), .IN6(na215_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na672_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x85y66     80'h00_0018_00_0010_0666_00FA
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a677_1 ( .OUT(na677_1), .IN1(na221_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na675_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y38     80'h00_0078_00_0020_0C66_FAFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a679_1 ( .OUT(na679_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na41_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na673_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a679_4 ( .OUT(na679_2), .COUTY1(na679_4), .IN1(1'b1), .IN2(na46_1), .IN3(1'b1), .IN4(1'b1), .IN5(na41_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na673_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x85y39     80'h00_0078_00_0020_0C66_AFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a681_1 ( .OUT(na681_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na50_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na679_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a681_4 ( .OUT(na681_2), .COUTY1(na681_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na54_1), .IN5(1'b1), .IN6(1'b1), .IN7(na50_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na679_4), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0018_0018_0014)) 
           _a685 ( .GLB0(na685_1), .GLB1(na685_2), .GLB2(na685_3), .GLB3(_d0), .CLK_FB0(_d1), .CLK_FB1(_d2), .CLK_FB2(_d3), .CLK_FB3(_d4),
                   .CLK0_0(na895_6), .CLK0_90(na895_5), .CLK0_180(na895_4), .CLK0_270(na895_3), .CLK0_BYP(1'b0), .CLK1_0(1'b0), .CLK1_90(1'b0),
                   .CLK1_180(1'b0), .CLK1_270(1'b0), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0), .CLK2_270(1'b0),
                   .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0), .USR_GLB0(1'b0),
                   .USR_GLB1(na897_9), .USR_GLB2(na904_9), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0), .USR_FB3(1'b0) );
// C_AND/D//AND/D      x96y39     80'h00_FA00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a703_1 ( .OUT(na703_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na272_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a703_2 ( .OUT(na703_1), .CLK(na685_1), .EN(na260_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na703_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a703_4 ( .OUT(na703_2_i), .IN1(na278_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a703_5 ( .OUT(na703_2), .CLK(na685_1), .EN(na260_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na703_2_i) );
// C_AND/D//AND/D      x96y42     80'h00_FA00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a704_1 ( .OUT(na704_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na274_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a704_2 ( .OUT(na704_1), .CLK(na685_1), .EN(na260_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na704_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a704_4 ( .OUT(na704_2_i), .IN1(na276_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a704_5 ( .OUT(na704_2), .CLK(na685_1), .EN(na260_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na704_2_i) );
// C_///AND/D      x95y29     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a707_4 ( .OUT(na707_2_i), .IN1(na280_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a707_5 ( .OUT(na707_2), .CLK(na685_1), .EN(na260_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na707_2_i) );
// C_AND/D///      x92y29     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a708_1 ( .OUT(na708_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na282_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a708_2 ( .OUT(na708_1), .CLK(na685_1), .EN(na260_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na708_1_i) );
// C_AND/D///      x94y30     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a709_1 ( .OUT(na709_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na283_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a709_2 ( .OUT(na709_1), .CLK(na685_1), .EN(na260_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na709_1_i) );
// C_AND/D///      x87y30     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a710_1 ( .OUT(na710_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na284_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a710_2 ( .OUT(na710_1), .CLK(na685_1), .EN(na260_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na710_1_i) );
// C_///AND/D      x88y33     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a717_4 ( .OUT(na717_2_i), .IN1(1'b1), .IN2(na468_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a717_5 ( .OUT(na717_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na717_2_i) );
// C_AND/D///      x88y31     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a719_1 ( .OUT(na719_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na490_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a719_2 ( .OUT(na719_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na719_1_i) );
// C_///AND/D      x90y35     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a721_4 ( .OUT(na721_2_i), .IN1(1'b1), .IN2(na512_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a721_5 ( .OUT(na721_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na721_2_i) );
// C_///AND/D      x90y34     80'h00_EE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a723_4 ( .OUT(na723_2_i), .IN1(na528_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a723_5 ( .OUT(na723_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na723_2_i) );
// C_///AND/D      x91y41     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a725_4 ( .OUT(na725_2_i), .IN1(1'b1), .IN2(na530_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a725_5 ( .OUT(na725_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na725_2_i) );
// C_AND/D///      x92y42     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a727_1 ( .OUT(na727_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na469_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a727_2 ( .OUT(na727_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na727_1_i) );
// C_///AND/D      x94y41     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a729_4 ( .OUT(na729_2_i), .IN1(1'b1), .IN2(na471_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a729_5 ( .OUT(na729_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na729_2_i) );
// C_AND/D///      x92y43     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a731_1 ( .OUT(na731_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na473_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a731_2 ( .OUT(na731_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na731_1_i) );
// C_AND/D///      x80y39     80'h00_EE00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a733_1 ( .OUT(na733_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na475_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a733_2 ( .OUT(na733_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na733_1_i) );
// C_AND/D///      x93y39     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a735_1 ( .OUT(na735_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na477_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a735_2 ( .OUT(na735_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na735_1_i) );
// C_///AND/D      x91y44     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a737_4 ( .OUT(na737_2_i), .IN1(1'b1), .IN2(na480_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a737_5 ( .OUT(na737_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na737_2_i) );
// C_AND/D///      x93y45     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a739_1 ( .OUT(na739_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na482_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a739_2 ( .OUT(na739_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na739_1_i) );
// C_///AND/D      x94y43     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a741_4 ( .OUT(na741_2_i), .IN1(1'b1), .IN2(na484_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a741_5 ( .OUT(na741_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na741_2_i) );
// C_///AND/D      x94y49     80'h00_EE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a743_4 ( .OUT(na743_2_i), .IN1(na486_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a743_5 ( .OUT(na743_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na743_2_i) );
// C_///AND/D      x90y51     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a745_4 ( .OUT(na745_2_i), .IN1(1'b1), .IN2(na488_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a745_5 ( .OUT(na745_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na745_2_i) );
// C_AND/D///      x90y51     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a747_1 ( .OUT(na747_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na491_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a747_2 ( .OUT(na747_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na747_1_i) );
// C_AND/D///      x92y53     80'h00_EE00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a749_1 ( .OUT(na749_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na493_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a749_2 ( .OUT(na749_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na749_1_i) );
// C_AND/D///      x94y52     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a751_1 ( .OUT(na751_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na495_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a751_2 ( .OUT(na751_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na751_1_i) );
// C_///AND/D      x92y51     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a753_4 ( .OUT(na753_2_i), .IN1(1'b1), .IN2(na497_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a753_5 ( .OUT(na753_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na753_2_i) );
// C_///AND/D      x90y55     80'h00_EE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a755_4 ( .OUT(na755_2_i), .IN1(na499_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a755_5 ( .OUT(na755_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na755_2_i) );
// C_///AND/D      x92y55     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a757_4 ( .OUT(na757_2_i), .IN1(1'b1), .IN2(na502_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a757_5 ( .OUT(na757_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na757_2_i) );
// C_AND/D///      x92y56     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a759_1 ( .OUT(na759_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na504_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a759_2 ( .OUT(na759_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na759_1_i) );
// C_///AND/D      x91y56     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a761_4 ( .OUT(na761_2_i), .IN1(1'b1), .IN2(na506_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a761_5 ( .OUT(na761_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na761_2_i) );
// C_AND/D///      x92y54     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a763_1 ( .OUT(na763_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na508_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a763_2 ( .OUT(na763_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na763_1_i) );
// C_AND/D///      x92y55     80'h00_EE00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a765_1 ( .OUT(na765_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na510_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a765_2 ( .OUT(na765_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na765_1_i) );
// C_AND/D///      x91y61     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a767_1 ( .OUT(na767_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na513_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a767_2 ( .OUT(na767_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na767_1_i) );
// C_///AND/D      x90y62     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a769_4 ( .OUT(na769_2_i), .IN1(1'b1), .IN2(na515_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a769_5 ( .OUT(na769_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na769_2_i) );
// C_AND/D///      x90y63     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a771_1 ( .OUT(na771_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na517_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a771_2 ( .OUT(na771_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na771_1_i) );
// C_///AND/D      x79y56     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a773_4 ( .OUT(na773_2_i), .IN1(1'b1), .IN2(na519_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a773_5 ( .OUT(na773_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na773_2_i) );
// C_///AND/D      x80y57     80'h00_EE00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a775_4 ( .OUT(na775_2_i), .IN1(na521_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a775_5 ( .OUT(na775_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na775_2_i) );
// C_///AND/D      x80y55     80'h00_EE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a777_4 ( .OUT(na777_2_i), .IN1(1'b1), .IN2(na524_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a777_5 ( .OUT(na777_2), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na777_2_i) );
// C_AND/D///      x80y55     80'h00_EE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a779_1 ( .OUT(na779_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na526_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a779_2 ( .OUT(na779_1), .CLK(na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na779_1_i) );
// C_AND/D//AND/D      x80y66     80'h00_ED00_80_0000_0C88_3FCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a780_1 ( .OUT(na780_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na780_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a780_2 ( .OUT(na780_1), .CLK(~na685_3), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na780_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a780_4 ( .OUT(na780_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na780_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a780_5 ( .OUT(na780_2), .CLK(~na685_3), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na780_2_i) );
// C_///AND/D      x77y55     80'h00_ED00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a782_4 ( .OUT(na782_2_i), .IN1(na463_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a782_5 ( .OUT(na782_2), .CLK(~na685_3), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na782_2_i) );
// C_AND/D///      x82y66     80'h00_ED00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a784_1 ( .OUT(na784_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na465_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a784_2 ( .OUT(na784_1), .CLK(~na685_3), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na784_1_i) );
// C_AND/D///      x79y65     80'h00_ED00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a788_1 ( .OUT(na788_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na685_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a788_2 ( .OUT(na788_1), .CLK(~na685_3), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na788_1_i) );
// C_AND/D///      x79y30     80'h00_EE00_00_0000_0C88_F3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a789_1 ( .OUT(na789_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na789_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a789_2 ( .OUT(na789_1), .CLK(na685_1), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na789_1_i) );
// C_///AND/D      x80y63     80'h00_EE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a791_4 ( .OUT(na791_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na460_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a791_5 ( .OUT(na791_2), .CLK(na685_1), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na791_2_i) );
// C_AND/D//AND/D      x88y29     80'h00_FE00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a857_1 ( .OUT(na857_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na857_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a857_2 ( .OUT(na857_1), .CLK(na685_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na857_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a857_4 ( .OUT(na857_2_i), .IN1(na894_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a857_5 ( .OUT(na857_2), .CLK(na685_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na857_2_i) );
// C_MX4a////      x79y51     80'h00_0018_00_0040_0C0A_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a869_1 ( .OUT(na869_1), .IN1(1'b0), .IN2(na1271_2), .IN3(1'b0), .IN4(na958_1), .IN5(na896_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1255_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x79y50     80'h00_0018_00_0040_0C05_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a870_1 ( .OUT(na870_1), .IN1(na1272_2), .IN2(1'b0), .IN3(na965_1), .IN4(1'b0), .IN5(~na896_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1255_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x80y49     80'h00_0018_00_0040_0C0A_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a871_1 ( .OUT(na871_1), .IN1(1'b0), .IN2(na1273_2), .IN3(1'b0), .IN4(na970_1), .IN5(na896_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1255_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x78y48     80'h00_0018_00_0040_0C05_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a872_1 ( .OUT(na872_1), .IN1(na1274_2), .IN2(1'b0), .IN3(na975_1), .IN4(1'b0), .IN5(~na896_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1255_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x80y54     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a873_1 ( .OUT(na873_1), .IN1(na782_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1256_2), .IN5(na869_1), .IN6(na870_1), .IN7(na871_1),
                     .IN8(na872_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x79y47     80'h00_0018_00_0040_0C0A_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a874_1 ( .OUT(na874_1), .IN1(1'b0), .IN2(na1275_2), .IN3(1'b0), .IN4(na978_1), .IN5(na896_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1255_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x79y46     80'h00_0018_00_0040_0C05_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a875_1 ( .OUT(na875_1), .IN1(na1277_2), .IN2(1'b0), .IN3(na986_1), .IN4(1'b0), .IN5(~na896_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1255_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x80y45     80'h00_0018_00_0040_0C0A_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a876_1 ( .OUT(na876_1), .IN1(1'b0), .IN2(na1278_2), .IN3(1'b0), .IN4(na991_1), .IN5(na896_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1255_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x78y44     80'h00_0018_00_0040_0C05_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a877_1 ( .OUT(na877_1), .IN1(na1279_2), .IN2(1'b0), .IN3(na993_1), .IN4(1'b0), .IN5(~na896_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1255_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x79y54     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a878_1 ( .OUT(na878_1), .IN1(na782_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1256_2), .IN5(na874_1), .IN6(na875_1), .IN7(na876_1),
                     .IN8(na877_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_04_05_00_02_80_01_00_00_00_03_03_00_00_00_33_03_13_33_00_00),
             .INIT_00(320'h0000000000095e1092c7000000000008faa08c8b00000000000896a0864700000000000832307fff),
             .INIT_01(320'h00000000000ae100ab1e00000000000a8260a52700000000000a22309f19000000000009c0a098f8),
             .INIT_02(320'h00000000000c47a0c1cd00000000000bf160bc5500000000000b98c0b6b900000000000b3de0b0fb),
             .INIT_03(320'h00000000000d8420d5f400000000000d39a0d13200000000000cebf0cc3f00000000000c9b30c71c),
             .INIT_04(320'h00000000000e8a50e6ce00000000000e4e70e2f100000000000e0eb0ded600000000000dcb30da81),
             .INIT_05(320'h00000000000f5030f3b400000000000f2540f0e100000000000ef5e0edc900000000000ec230ea6c),
             .INIT_06(320'h00000000000fce20fc2800000000000fb5c0fa7c00000000000f9890f88300000000000f76b0f640),
             .INIT_07(320'h00000000000fff50ffd700000000000ffa60ff6100000000000ff080fe9c00000000000fe1c0fd89),
             .INIT_08(320'h00000000000fe1c0fe9c00000000000ff080ff6100000000000ffa60ffd700000000000fff50ffff),
             .INIT_09(320'h00000000000f76b0f88300000000000f9890fa7c00000000000fb5c0fc2800000000000fce20fd89),
             .INIT_0A(320'h00000000000ec230edc900000000000ef5e0f0e100000000000f2540f3b400000000000f5030f640),
             .INIT_0B(320'h00000000000dcb30ded600000000000e0eb0e2f100000000000e4e70e6ce00000000000e8a50ea6c),
             .INIT_0C(320'h00000000000c9b30cc3f00000000000cebf0d13200000000000d39a0d5f400000000000d8420da81),
             .INIT_0D(320'h00000000000b3de0b6b900000000000b98c0bc5500000000000bf160c1cd00000000000c47a0c71c),
             .INIT_0E(320'h000000000009c0a09f1900000000000a2230a52700000000000a8260ab1e00000000000ae100b0fb),
             .INIT_0F(320'h0000000000083230864700000000000896a08c8b000000000008faa092c70000000000095e1098f8),
             .INIT_10(320'h000000000006a1d06d3700000000000705407373000000000007694079b7000000000007cdb07fff),
             .INIT_11(320'h0000000000051ee054e00000000000057d805ad7000000000005ddb060e50000000000063f406706),
             .INIT_12(320'h000000000003b8403e310000000000040e8043a900000000000467204945000000000004c2004f03),
             .INIT_13(320'h0000000000027bc02a0a000000000002c6402ecc00000000000313f033bf00000000000364b038e2),
             .INIT_14(320'h00000000000175901930000000000001b1701d0d000000000001f130212800000000000234b0257d),
             .INIT_15(320'h000000000000afb00c4a000000000000daa00f1d0000000000010a0012350000000000013db01592),
             .INIT_16(320'h00000000000031c003d60000000000004a2005820000000000006750077b000000000000893009be),
             .INIT_17(320'h000000000000009000270000000000000580009d0000000000000f6001620000000000001e200275),
             .INIT_18(320'h0000000000001e2001620000000000000f60009d0000000000000580002700000000000000900000),
             .INIT_19(320'h0000000000008930077b000000000000675005820000000000004a2003d600000000000031c00275),
             .INIT_1A(320'h0000000000013db012350000000000010a000f1d000000000000daa00c4a000000000000afb009be),
             .INIT_1B(320'h00000000000234b02128000000000001f1301d0d000000000001b170193000000000000175901592),
             .INIT_1C(320'h00000000000364b033bf00000000000313f02ecc000000000002c6402a0a0000000000027bc0257d),
             .INIT_1D(320'h000000000004c2004945000000000004672043a90000000000040e803e31000000000003b84038e2),
             .INIT_1E(320'h0000000000063f4060e5000000000005ddb05ad70000000000057d8054e00000000000051ee04f03),
             .INIT_1F(320'h000000000007cdb079b70000000000076940737300000000000705406d37000000000006a1d06706),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a879 ( .DOA({_d5, _d6, _d7, _d8, _d9, _d10, _d11, _d12, _d13, _d14, _d15, _d16, _d17, _d18, _d19, _d20, _d21, _d22, _d23,
                  _d24, _d25, _d26, _d27, _d28, na879_25, na879_26, na879_27, na879_28, na879_29, na879_30, na879_31, na879_32, na879_33,
                  na879_34, na879_35, na879_36, na879_37, na879_38, na879_39, na879_40}),
                   .DOAX({_d29, _d30, _d31, _d32, _d33, _d34, _d35, _d36, _d37, _d38, _d39, _d40, _d41, _d42, _d43, _d44, _d45, _d46,
                  _d47, _d48, _d49, _d50, _d51, _d52, _d53, _d54, _d55, _d56, _d57, _d58, _d59, _d60, _d61, _d62, _d63, _d64, _d65,
                  _d66, _d67, _d68}),
                   .DOB({_d69, _d70, _d71, _d72, _d73, _d74, _d75, _d76, _d77, _d78, _d79, _d80, _d81, _d82, _d83, _d84, _d85, _d86,
                  _d87, _d88, _d89, _d90, _d91, _d92, _d93, _d94, _d95, _d96, _d97, _d98, _d99, _d100, _d101, _d102, _d103, _d104,
                  _d105, _d106, _d107, _d108}),
                   .DOBX({_d109, _d110, _d111, _d112, _d113, _d114, _d115, _d116, _d117, _d118, _d119, _d120, _d121, _d122, _d123,
                  _d124, _d125, _d126, _d127, _d128, _d129, _d130, _d131, _d132, _d133, _d134, _d135, _d136, _d137, _d138, _d139, _d140,
                  _d141, _d142, _d143, _d144, _d145, _d146, _d147, _d148}),
                   .ECC1B_ERRA({_d149, _d150, _d151, _d152}),
                   .ECC1B_ERRB({_d153, _d154, _d155, _d156}),
                   .ECC2B_ERRA({_d157, _d158, _d159, _d160}),
                   .ECC2B_ERRB({_d161, _d162, _d163, _d164}),
                   .FORW_CAS_WRAO(_d165), .FORW_CAS_WRBO(_d166), .FORW_CAS_BMAO(_d167), .FORW_CAS_BMBO(_d168), .FORW_CAS_RDAO(_d169),
                   .FORW_CAS_RDBO(_d170), .FORW_UADDRAO({_d171, _d172, _d173, _d174, _d175, _d176, _d177, _d178, _d179, _d180, _d181,
                  _d182, _d183, _d184, _d185, _d186}),
                   .FORW_LADDRAO({_d187, _d188, _d189, _d190, _d191, _d192, _d193, _d194, _d195, _d196, _d197, _d198, _d199, _d200,
                  _d201, _d202}),
                   .FORW_UADDRBO({_d203, _d204, _d205, _d206, _d207, _d208, _d209, _d210, _d211, _d212, _d213, _d214, _d215, _d216,
                  _d217, _d218}),
                   .FORW_LADDRBO({_d219, _d220, _d221, _d222, _d223, _d224, _d225, _d226, _d227, _d228, _d229, _d230, _d231, _d232,
                  _d233, _d234}),
                   .FORW_UA0CLKO(_d235), .FORW_UA0ENO(_d236), .FORW_UA0WEO(_d237), .FORW_LA0CLKO(_d238), .FORW_LA0ENO(_d239), .FORW_LA0WEO(_d240),
                   .FORW_UA1CLKO(_d241), .FORW_UA1ENO(_d242), .FORW_UA1WEO(_d243), .FORW_LA1CLKO(_d244), .FORW_LA1ENO(_d245), .FORW_LA1WEO(_d246),
                   .FORW_UB0CLKO(_d247), .FORW_UB0ENO(_d248), .FORW_UB0WEO(_d249), .FORW_LB0CLKO(_d250), .FORW_LB0ENO(_d251), .FORW_LB0WEO(_d252),
                   .FORW_UB1CLKO(_d253), .FORW_UB1ENO(_d254), .FORW_UB1WEO(_d255), .FORW_LB1CLKO(_d256), .FORW_LB1ENO(_d257), .FORW_LB1WEO(_d258),
                   .CLOCKA({_d259, _d260, _d261, _d262}),
                   .CLOCKB({_d263, _d264, _d265, _d266}),
                   .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .CLKB({1'b1, 1'b1, 1'b1, na907_9}),
                   .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .GLWEA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0({na908_10, na909_9, na910_10, na911_9, na915_10, na917_9, na918_10, na922_9, na923_10, na928_9, na929_10,
                  na932_9, na934_10, na935_9, na937_10, na940_9}),
                   .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na943_9, 1'b1, na946_9, na947_10, na948_9, na952_10,
                  na953_9}),
                   .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .CLOCK1(1'b1), .CLOCK2(na685_2), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                   .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                   .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                   .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                   .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a880 ( .Y(na880_1), .I(arst_n) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a881 ( .O(bck), .A(na1204_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a882 ( .Y(na882_1), .I(clk) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a883 ( .O(clk_check), .A(na1205_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a884 ( .O(din), .A(na1206_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a885 ( .O(led[0]), .A(na1207_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a886 ( .O(led[1]), .A(na1208_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a887 ( .O(led[2]), .A(na1209_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a888 ( .O(led[3]), .A(na1210_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a889 ( .O(led[4]), .A(na1211_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a890 ( .O(led[5]), .A(na1212_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a891 ( .O(led[6]), .A(na1213_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a892 ( .O(led[7]), .A(na1214_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a893 ( .O(lrck), .A(na1215_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a894 ( .Y(na894_1), .I(uart_rx_serial) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_05_08_0C_20_82)) 
           _a895 ( .USR_PLL_LOCKED_STDY(_d267), .USR_PLL_LOCKED(_d268), .CLK270(na895_3), .CLK180(na895_4), .CLK90(na895_5), .CLK0(na895_6),
                   .CLK_REF_OUT(_d269), .CLK_REF(na906_1), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
// C_///AND/D      x79y45     80'h00_ED00_80_0000_0C08_FFFF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a896_4 ( .OUT(na896_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a896_5 ( .OUT(na896_2), .CLK(~na685_2), .EN(1'b1), .SR(na880_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na896_2_i) );
// C_AND////      x1y127     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a897_1 ( .OUT(na897_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na467_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a897_6 ( .RAM_O1(na897_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na897_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x85y34     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a898_2 ( .OUT(na898_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a898_6 ( .COUTY1(na898_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na898_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x81y35     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a899_1 ( .OUT(na899_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na406_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x82y37     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a900_1 ( .OUT(na900_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na629_1), .IN6(na1222_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x93y38     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a901_1 ( .OUT(na901_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0), .CINX(1'b0),
                     .CINY1(na322_4), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y36     80'h00_0078_00_0000_0CEE_5555
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a902_1 ( .OUT(na902_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na406_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a902_4 ( .OUT(na902_2), .IN1(~na629_2), .IN2(1'b0), .IN3(~na1220_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y35     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a903_4 ( .OUT(na903_2), .IN1(1'b1), .IN2(na22_2), .IN3(na343_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x1y126     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a904_1 ( .OUT(na904_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na791_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a904_6 ( .RAM_O1(na904_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na904_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x91y42     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a905_4 ( .OUT(na905_2), .IN1(1'b1), .IN2(na22_1), .IN3(na566_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a906 ( .PCLK0(na906_1), .PCLK1(_d270), .PCLK2(_d271), .PCLK3(_d272), .CLK0(na882_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0),
                   .SER_CLK(1'b0), .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_AND////      x67y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a907_1 ( .OUT(na907_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a907_6 ( .RAM_O1(na907_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na907_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a908_4 ( .OUT(na908_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a908_6 ( .RAM_O2(na908_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na908_2), .COMP_OUT(1'b0) );
// C_AND////      x60y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a909_1 ( .OUT(na909_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a909_6 ( .RAM_O1(na909_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na909_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y39     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a910_4 ( .OUT(na910_2), .IN1(1'b1), .IN2(1'b1), .IN3(na779_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a910_6 ( .RAM_O2(na910_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na910_2), .COMP_OUT(1'b0) );
// C_AND////      x60y39     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a911_1 ( .OUT(na911_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na526_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a911_6 ( .RAM_O1(na911_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na911_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x84y31     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a912_1 ( .OUT(na912_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0), .CINX(1'b0),
                     .CINY1(na552_4), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x83y37     80'h00_0078_00_0000_0CEE_5555
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a913_1 ( .OUT(na913_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na450_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a913_4 ( .OUT(na913_2), .IN1(~na673_1), .IN2(1'b0), .IN3(~na1220_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x82y37     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a914_4 ( .OUT(na914_2), .IN1(1'b1), .IN2(na22_2), .IN3(1'b1), .IN4(na365_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y38     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a915_4 ( .OUT(na915_2), .IN1(1'b1), .IN2(1'b1), .IN3(na777_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a915_6 ( .RAM_O2(na915_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na915_2), .COMP_OUT(1'b0) );
// C_AND////      x83y36     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a916_1 ( .OUT(na916_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na588_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y38     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a917_1 ( .OUT(na917_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na524_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a917_6 ( .RAM_O1(na917_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na917_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y37     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a918_4 ( .OUT(na918_2), .IN1(1'b1), .IN2(1'b1), .IN3(na775_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a918_6 ( .RAM_O2(na918_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na918_2), .COMP_OUT(1'b0) );
// C_AND////      x94y42     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a919_1 ( .OUT(na919_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na610_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y38     80'h00_0078_00_0000_0CEE_5555
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a920_1 ( .OUT(na920_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na673_2), .IN6(1'b0), .IN7(~na1220_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a920_4 ( .OUT(na920_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na450_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x81y41     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a921_1 ( .OUT(na921_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(na387_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y37     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a922_1 ( .OUT(na922_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na521_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a922_6 ( .RAM_O1(na922_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na922_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y36     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a923_4 ( .OUT(na923_2), .IN1(1'b1), .IN2(na773_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a923_6 ( .RAM_O2(na923_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na923_2), .COMP_OUT(1'b0) );
// C_///AND/      x81y41     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a924_4 ( .OUT(na924_2), .IN1(1'b1), .IN2(na22_2), .IN3(na387_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x81y44     80'h00_0078_00_0000_0CEE_0735
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a925_1 ( .OUT(na925_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_1), .IN6(~na679_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a925_4 ( .OUT(na925_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na456_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y40     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a926_4 ( .OUT(na926_2), .IN1(1'b1), .IN2(na22_1), .IN3(na610_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x81y46     80'h00_0078_00_0000_0C88_CCF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a927_1 ( .OUT(na927_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na615_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a927_4 ( .OUT(na927_2), .IN1(na10_1), .IN2(na679_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a928_1 ( .OUT(na928_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a928_6 ( .RAM_O1(na928_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na928_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x60y35     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a929_4 ( .OUT(na929_2), .IN1(1'b1), .IN2(na519_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a929_6 ( .RAM_O2(na929_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na929_2), .COMP_OUT(1'b0) );
// C_OR///OR/      x91y39     80'h00_0078_00_0000_0CEE_5555
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a930_1 ( .OUT(na930_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na458_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a930_4 ( .OUT(na930_2), .IN1(~na681_1), .IN2(1'b0), .IN3(~na1220_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y44     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a931_1 ( .OUT(na931_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na615_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y35     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a932_1 ( .OUT(na932_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a932_6 ( .RAM_O1(na932_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na932_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x83y40     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a933_4 ( .OUT(na933_2), .IN1(1'b1), .IN2(na22_2), .IN3(1'b1), .IN4(na392_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y34     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a934_4 ( .OUT(na934_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a934_6 ( .RAM_O2(na934_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na934_2), .COMP_OUT(1'b0) );
// C_AND////      x60y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a935_1 ( .OUT(na935_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a935_6 ( .RAM_O1(na935_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na935_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x81y47     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a936_1 ( .OUT(na936_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na681_2), .IN6(na1222_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a937_4 ( .OUT(na937_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a937_6 ( .RAM_O2(na937_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na937_2), .COMP_OUT(1'b0) );
// C_OR///OR/      x81y38     80'h00_0078_00_0000_0CEE_5355
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a938_1 ( .OUT(na938_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(~na394_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a938_4 ( .OUT(na938_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na458_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x96y47     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a939_4 ( .OUT(na939_2), .IN1(1'b1), .IN2(na22_1), .IN3(na617_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a940_1 ( .OUT(na940_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a940_6 ( .RAM_O1(na940_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na940_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR///OR/      x82y39     80'h00_0078_00_0000_0CEE_5335
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a941_1 ( .OUT(na941_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(~na394_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a941_4 ( .OUT(na941_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na397_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x83y40     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a942_1 ( .OUT(na942_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na617_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a943_1 ( .OUT(na943_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a943_6 ( .RAM_O1(na943_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na943_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x81y47     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a944_4 ( .OUT(na944_2), .IN1(na10_1), .IN2(na620_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x90y40     80'h00_0078_00_0000_0C88_CCF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a945_1 ( .OUT(na945_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na557_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a945_4 ( .OUT(na945_2), .IN1(na10_1), .IN2(na620_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x69y35     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a946_1 ( .OUT(na946_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a946_6 ( .RAM_O1(na946_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na946_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x69y34     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a947_4 ( .OUT(na947_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a947_6 ( .RAM_O2(na947_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na947_2), .COMP_OUT(1'b0) );
// C_AND////      x69y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a948_1 ( .OUT(na948_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a948_6 ( .RAM_O1(na948_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na948_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x92y47     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a949_1 ( .OUT(na949_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na557_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x80y40     80'h00_0078_00_0000_0CEE_5533
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a950_1 ( .OUT(na950_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na399_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a950_4 ( .OUT(na950_2), .IN1(1'b0), .IN2(~na22_2), .IN3(1'b0), .IN4(~na334_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y49     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a951_4 ( .OUT(na951_2), .IN1(na622_1), .IN2(na1222_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a952_4 ( .OUT(na952_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a952_6 ( .RAM_O2(na952_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na952_2), .COMP_OUT(1'b0) );
// C_AND////      x69y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a953_1 ( .OUT(na953_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a953_6 ( .RAM_O1(na953_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na953_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x79y40     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a954_4 ( .OUT(na954_2), .IN1(1'b1), .IN2(na22_2), .IN3(na336_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y41     80'h00_0078_00_0000_0CEE_5555
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a955_1 ( .OUT(na955_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na399_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a955_4 ( .OUT(na955_2), .IN1(~na622_2), .IN2(1'b0), .IN3(~na1220_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y43     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a956_1 ( .OUT(na956_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na559_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x64y40     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a957_5 ( .OUT(na957_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_25), .CP_O(1'b0) );
// C_/RAM_I1///      x64y40     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a958_2 ( .OUT(na958_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_26), .CP_O(1'b0) );
// C_///AND/      x92y44     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a959_4 ( .OUT(na959_2), .IN1(1'b1), .IN2(na22_1), .IN3(na559_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x81y42     80'h00_0078_00_0000_0CEE_3507
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a960_1 ( .OUT(na960_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na401_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a960_4 ( .OUT(na960_2), .IN1(~na10_1), .IN2(~na624_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x78y43     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a961_1 ( .OUT(na961_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(na336_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x64y39     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a962_5 ( .OUT(na962_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_27), .CP_O(1'b0) );
// C_OR///OR/      x81y43     80'h00_0078_00_0000_0CEE_0735
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a963_1 ( .OUT(na963_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_1), .IN6(~na624_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a963_4 ( .OUT(na963_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na401_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y47     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a964_4 ( .OUT(na964_2), .IN1(1'b1), .IN2(na22_1), .IN3(1'b1), .IN4(na561_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x64y39     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a965_2 ( .OUT(na965_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_28), .CP_O(1'b0) );
// C_AND////      x90y39     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a966_1 ( .OUT(na966_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(1'b1), .IN8(na338_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x64y38     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a967_5 ( .OUT(na967_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_29), .CP_O(1'b0) );
// C_OR///OR/      x82y44     80'h00_0078_00_0000_0CEE_3355
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a968_1 ( .OUT(na968_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(1'b0), .IN8(~na338_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a968_4 ( .OUT(na968_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na403_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y46     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a969_1 ( .OUT(na969_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na561_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x64y38     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a970_2 ( .OUT(na970_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_30), .CP_O(1'b0) );
// C_AND////      x81y49     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a971_1 ( .OUT(na971_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na626_1), .IN6(na1222_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x64y37     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a972_5 ( .OUT(na972_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_31), .CP_O(1'b0) );
// C_OR///OR/      x80y44     80'h00_0078_00_0000_0CEE_5555
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a973_1 ( .OUT(na973_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na403_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a973_4 ( .OUT(na973_2), .IN1(~na626_2), .IN2(1'b0), .IN3(~na1220_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x79y41     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a974_4 ( .OUT(na974_2), .IN1(1'b1), .IN2(na22_2), .IN3(na340_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x64y37     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a975_2 ( .OUT(na975_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_32), .CP_O(1'b0) );
// C_AND////      x94y43     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a976_1 ( .OUT(na976_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na563_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x64y36     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a977_5 ( .OUT(na977_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_33), .CP_O(1'b0) );
// C_/RAM_I1///      x64y36     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a978_2 ( .OUT(na978_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_34), .CP_O(1'b0) );
// C_///AND/      x78y40     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a979_4 ( .OUT(na979_2), .IN1(1'b1), .IN2(na22_2), .IN3(na340_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y45     80'h00_0078_00_0000_0CEE_3507
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a980_1 ( .OUT(na980_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na405_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a980_4 ( .OUT(na980_2), .IN1(~na10_1), .IN2(~na628_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y45     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a981_1 ( .OUT(na981_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na563_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x92y48     80'h00_0078_00_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a982_1 ( .OUT(na982_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(1'b1), .IN8(na342_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a982_4 ( .OUT(na982_2), .IN1(1'b1), .IN2(na22_1), .IN3(1'b1), .IN4(na565_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x64y35     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a983_5 ( .OUT(na983_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_35), .CP_O(1'b0) );
// C_///OR/      x85y34     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a984_4 ( .OUT(na984_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na405_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x83y34     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a985_4 ( .OUT(na985_2), .IN1(na10_1), .IN2(na628_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x64y35     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a986_2 ( .OUT(na986_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_36), .CP_O(1'b0) );
// C_OR///OR/      x82y47     80'h00_0078_00_0000_0CEE_3355
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a987_1 ( .OUT(na987_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(1'b0), .IN8(~na342_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a987_4 ( .OUT(na987_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na408_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y46     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a988_1 ( .OUT(na988_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na565_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x64y34     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a989_5 ( .OUT(na989_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_37), .CP_O(1'b0) );
// C_///AND/      x80y48     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a990_4 ( .OUT(na990_2), .IN1(na631_1), .IN2(na1222_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x64y34     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a991_2 ( .OUT(na991_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_38), .CP_O(1'b0) );
// C_////RAM_I2      x64y33     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a992_5 ( .OUT(na992_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_39), .CP_O(1'b0) );
// C_/RAM_I1///      x64y33     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a993_2 ( .OUT(na993_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na879_40), .CP_O(1'b0) );
// C_OR///OR/      x82y46     80'h00_0078_00_0000_0CEE_3553
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a995_1 ( .OUT(na995_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na410_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a995_4 ( .OUT(na995_2), .IN1(1'b0), .IN2(~na22_2), .IN3(~na345_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y51     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a996_1 ( .OUT(na996_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na10_1), .IN6(na633_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y46     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a998_4 ( .OUT(na998_2), .IN1(1'b1), .IN2(na22_1), .IN3(na568_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x80y47     80'h00_0078_00_0000_0CEE_3507
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1000_1 ( .OUT(na1000_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na410_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1000_4 ( .OUT(na1000_2), .IN1(~na10_1), .IN2(~na633_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x80y52     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1001_1 ( .OUT(na1001_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(1'b1), .IN8(na347_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y44     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1003_4 ( .OUT(na1003_2), .IN1(1'b1), .IN2(na22_1), .IN3(1'b1), .IN4(na570_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y48     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1009_1 ( .OUT(na1009_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na635_2), .IN6(na1222_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y51     80'h00_0078_00_0000_0CEE_5355
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1010_1 ( .OUT(na1010_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(~na349_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1010_4 ( .OUT(na1010_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na412_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y50     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1011_4 ( .OUT(na1011_2), .IN1(1'b1), .IN2(na22_1), .IN3(na572_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x78y52     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1014_1 ( .OUT(na1014_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(na349_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x78y45     80'h00_0078_00_0000_0CEE_3507
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1015_1 ( .OUT(na1015_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na414_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1015_4 ( .OUT(na1015_2), .IN1(~na10_1), .IN2(~na637_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y48     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1016_4 ( .OUT(na1016_2), .IN1(1'b1), .IN2(na22_1), .IN3(na572_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x78y54     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1019_4 ( .OUT(na1019_2), .IN1(1'b1), .IN2(na22_2), .IN3(1'b1), .IN4(na351_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x81y53     80'h00_0078_00_0000_0CEE_0735
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1020_1 ( .OUT(na1020_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_1), .IN6(~na637_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1020_4 ( .OUT(na1020_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na414_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y48     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1021_1 ( .OUT(na1021_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na574_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x77y53     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1024_1 ( .OUT(na1024_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(1'b1), .IN8(na351_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y53     80'h00_0078_00_0000_0CEE_5555
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1025_1 ( .OUT(na1025_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na639_1), .IN6(1'b0), .IN7(~na1220_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1025_4 ( .OUT(na1025_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na416_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y54     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1026_1 ( .OUT(na1026_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na574_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y52     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1029_4 ( .OUT(na1029_2), .IN1(na639_2), .IN2(na1222_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y50     80'h00_0078_00_0000_0CEE_5355
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1030_1 ( .OUT(na1030_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(~na353_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1030_4 ( .OUT(na1030_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na416_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y50     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1031_1 ( .OUT(na1031_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na576_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x80y50     80'h00_0078_00_0000_0CEE_0735
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1033_1 ( .OUT(na1033_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_1), .IN6(~na642_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1033_4 ( .OUT(na1033_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na419_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y52     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1034_4 ( .OUT(na1034_2), .IN1(1'b1), .IN2(na22_1), .IN3(na576_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x80y53     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1036_1 ( .OUT(na1036_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(na353_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y52     80'h00_0078_00_0000_0CEE_3335
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1038_1 ( .OUT(na1038_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(1'b0), .IN8(~na356_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1038_4 ( .OUT(na1038_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na419_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y50     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1039_4 ( .OUT(na1039_2), .IN1(1'b1), .IN2(na22_1), .IN3(1'b1), .IN4(na579_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x82y55     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1041_1 ( .OUT(na1041_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na10_1), .IN6(na642_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y46     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1044_4 ( .OUT(na1044_2), .IN1(1'b1), .IN2(na22_1), .IN3(1'b1), .IN4(na579_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x81y51     80'h00_0078_00_0000_0CEE_5533
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1045_1 ( .OUT(na1045_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na421_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1045_4 ( .OUT(na1045_2), .IN1(1'b0), .IN2(~na22_2), .IN3(1'b0), .IN4(~na356_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y55     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1046_1 ( .OUT(na1046_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na644_1), .IN6(na1222_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x79y53     80'h00_0078_00_0000_0CEE_5555
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1048_1 ( .OUT(na1048_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na421_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1048_4 ( .OUT(na1048_2), .IN1(~na644_2), .IN2(1'b0), .IN3(~na1220_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y54     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1049_4 ( .OUT(na1049_2), .IN1(1'b1), .IN2(na22_2), .IN3(na358_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y53     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1051_1 ( .OUT(na1051_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na581_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x80y46     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1054_4 ( .OUT(na1054_2), .IN1(1'b1), .IN2(na22_2), .IN3(na358_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x81y54     80'h00_0078_00_0000_0CEE_0735
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1055_1 ( .OUT(na1055_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_1), .IN6(~na646_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1055_4 ( .OUT(na1055_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na423_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y48     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1056_4 ( .OUT(na1056_2), .IN1(1'b1), .IN2(na22_1), .IN3(na581_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x81y56     80'h00_0018_00_0000_0CEE_3500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1058_1 ( .OUT(na1058_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na423_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y56     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1059_4 ( .OUT(na1059_2), .IN1(na10_1), .IN2(na646_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x93y54     80'h00_0078_00_0000_0C88_CC88
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1060_1 ( .OUT(na1060_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na583_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1060_4 ( .OUT(na1060_2), .IN1(na9_2), .IN2(na7_1), .IN3(na425_1), .IN4(na1218_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x83y56     80'h00_0078_00_0000_0CEE_5555
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1063_1 ( .OUT(na1063_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na648_2), .IN6(1'b0), .IN7(~na1220_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1063_4 ( .OUT(na1063_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na425_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x79y45     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1064_1 ( .OUT(na1064_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(na362_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x96y55     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1066_4 ( .OUT(na1066_2), .IN1(1'b1), .IN2(na22_1), .IN3(na585_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x78y47     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1069_1 ( .OUT(na1069_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(na362_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x81y55     80'h00_0078_00_0000_0CEE_3507
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1070_1 ( .OUT(na1070_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na427_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1070_4 ( .OUT(na1070_2), .IN1(~na10_1), .IN2(~na650_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y50     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1071_1 ( .OUT(na1071_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na585_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y58     80'h00_0078_00_0000_0CEE_0735
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1073_1 ( .OUT(na1073_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_1), .IN6(~na650_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1073_4 ( .OUT(na1073_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na427_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y53     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1074_4 ( .OUT(na1074_2), .IN1(1'b1), .IN2(na22_1), .IN3(1'b1), .IN4(na587_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y59     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1076_1 ( .OUT(na1076_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(1'b1), .IN8(na364_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y56     80'h00_0078_00_0000_0CEE_3355
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1078_1 ( .OUT(na1078_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(1'b0), .IN8(~na364_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1078_4 ( .OUT(na1078_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na430_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y54     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1079_4 ( .OUT(na1079_2), .IN1(1'b1), .IN2(na22_1), .IN3(1'b1), .IN4(na587_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x82y57     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1081_1 ( .OUT(na1081_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na653_1), .IN6(na1222_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x81y58     80'h00_0078_00_0000_0CEE_5553
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1083_1 ( .OUT(na1083_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na430_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1083_4 ( .OUT(na1083_2), .IN1(1'b0), .IN2(~na22_2), .IN3(~na367_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x79y55     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1084_4 ( .OUT(na1084_2), .IN1(na653_2), .IN2(na1221_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y56     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1086_1 ( .OUT(na1086_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na590_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x92y57     80'h00_0078_00_0000_0CEE_3553
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1088_1 ( .OUT(na1088_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na432_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1088_4 ( .OUT(na1088_2), .IN1(1'b0), .IN2(~na22_2), .IN3(~na367_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x80y58     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1089_4 ( .OUT(na1089_2), .IN1(na10_1), .IN2(na655_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y56     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1091_4 ( .OUT(na1091_2), .IN1(1'b1), .IN2(na22_1), .IN3(na590_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x91y58     80'h00_0078_00_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1098_1 ( .OUT(na1098_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(na371_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1098_4 ( .OUT(na1098_2), .IN1(1'b1), .IN2(na22_1), .IN3(na594_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x80y56     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1100_4 ( .OUT(na1100_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na434_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x80y57     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1101_1 ( .OUT(na1101_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na657_2), .IN6(na1222_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x83y60     80'h00_0078_00_0000_0CEE_3507
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1103_1 ( .OUT(na1103_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na436_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1103_4 ( .OUT(na1103_2), .IN1(~na10_1), .IN2(~na659_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x82y55     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1104_4 ( .OUT(na1104_2), .IN1(1'b1), .IN2(na22_2), .IN3(na371_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y58     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1106_1 ( .OUT(na1106_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na594_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x82y59     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1109_4 ( .OUT(na1109_2), .IN1(na10_1), .IN2(na659_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y60     80'h00_0078_00_0000_0CEE_3335
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1110_1 ( .OUT(na1110_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(1'b0), .IN8(~na373_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1110_4 ( .OUT(na1110_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na436_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y56     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1111_1 ( .OUT(na1111_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na596_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y59     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1114_4 ( .OUT(na1114_2), .IN1(na661_1), .IN2(na1221_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x80y60     80'h00_0078_00_0000_0CEE_3355
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1115_1 ( .OUT(na1115_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(1'b0), .IN8(~na373_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1115_4 ( .OUT(na1115_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na438_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y50     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1116_1 ( .OUT(na1116_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na596_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y61     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1119_4 ( .OUT(na1119_2), .IN1(na661_2), .IN2(na1221_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x83y61     80'h00_0078_00_0000_0CEE_5355
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1120_1 ( .OUT(na1120_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(~na375_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1120_4 ( .OUT(na1120_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na438_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y58     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1121_1 ( .OUT(na1121_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na598_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x91y59     80'h00_0078_00_0000_0C88_F8AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1122_1 ( .OUT(na1122_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na10_1), .IN6(na664_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1122_4 ( .OUT(na1122_2), .IN1(1'b1), .IN2(na22_1), .IN3(na598_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x81y60     80'h00_0060_00_0000_0C0E_FF35
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1124_4 ( .OUT(na1124_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na441_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x80y58     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1125_1 ( .OUT(na1125_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(na375_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x94y59     80'h00_0078_00_0000_0C88_CCF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1126_1 ( .OUT(na1126_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na601_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1126_4 ( .OUT(na1126_2), .IN1(na10_1), .IN2(na664_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x81y61     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1130_4 ( .OUT(na1130_2), .IN1(na666_1), .IN2(na1221_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x81y62     80'h00_0078_00_0000_0CEE_3355
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1131_1 ( .OUT(na1131_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(1'b0), .IN8(~na378_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1131_4 ( .OUT(na1131_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na443_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y59     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1132_1 ( .OUT(na1132_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na601_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x92y63     80'h00_0078_00_0000_0CEE_5555
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1134_1 ( .OUT(na1134_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na443_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1134_4 ( .OUT(na1134_2), .IN1(~na666_2), .IN2(1'b0), .IN3(~na1220_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x78y56     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1135_4 ( .OUT(na1135_2), .IN1(1'b1), .IN2(na22_2), .IN3(na380_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y60     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1137_1 ( .OUT(na1137_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na603_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x82y59     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1140_1 ( .OUT(na1140_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na10_1), .IN6(na668_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y62     80'h00_0078_00_0000_0CEE_5335
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1141_1 ( .OUT(na1141_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(~na380_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1141_4 ( .OUT(na1141_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na445_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x93y61     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1142_1 ( .OUT(na1142_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na603_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x79y63     80'h00_0078_00_0000_0CEE_0735
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1144_1 ( .OUT(na1144_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_1), .IN6(~na668_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1144_4 ( .OUT(na1144_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na445_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y56     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1145_4 ( .OUT(na1145_2), .IN1(1'b1), .IN2(na22_1), .IN3(1'b1), .IN4(na605_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x81y60     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1147_1 ( .OUT(na1147_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_2), .IN7(1'b1), .IN8(na382_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x92y58     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1150_4 ( .OUT(na1150_2), .IN1(1'b1), .IN2(na22_1), .IN3(1'b1), .IN4(na605_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x84y65     80'h00_0078_00_0000_0CEE_5533
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1151_1 ( .OUT(na1151_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(~na447_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1151_4 ( .OUT(na1151_2), .IN1(1'b0), .IN2(~na22_2), .IN3(1'b0), .IN4(~na382_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x93y50     80'h00_0078_00_0000_0C88_AA18
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1152_1 ( .OUT(na1152_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na670_1), .IN6(1'b1), .IN7(na1220_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1152_4 ( .OUT(na1152_2), .IN1(na15_1), .IN2(na7_2), .IN3(~na703_2), .IN4(~na704_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y61     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1156_1 ( .OUT(na1156_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na607_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x83y64     80'h00_0078_00_0000_0CEE_3553
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1157_1 ( .OUT(na1157_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_2), .IN6(1'b0), .IN7(1'b0), .IN8(~na449_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1157_4 ( .OUT(na1157_2), .IN1(1'b0), .IN2(~na22_2), .IN3(~na384_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x91y61     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1158_4 ( .OUT(na1158_2), .IN1(na10_1), .IN2(na672_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x82y65     80'h00_0078_00_0000_0CEE_0735
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1160_1 ( .OUT(na1160_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na10_1), .IN6(~na672_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1160_4 ( .OUT(na1160_2), .IN1(~na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na449_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y62     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1161_1 ( .OUT(na1161_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(1'b1), .IN8(na609_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x78y58     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1163_4 ( .OUT(na1163_2), .IN1(1'b1), .IN2(na22_2), .IN3(1'b1), .IN4(na386_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x81y64     80'h00_0078_00_0000_0CEE_3355
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1165_1 ( .OUT(na1165_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na22_2), .IN7(1'b0), .IN8(~na386_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1165_4 ( .OUT(na1165_2), .IN1(~na10_2), .IN2(1'b0), .IN3(~na452_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y62     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1166_4 ( .OUT(na1166_2), .IN1(1'b1), .IN2(na22_1), .IN3(1'b1), .IN4(na609_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y63     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1168_1 ( .OUT(na1168_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na675_1), .IN6(na1221_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x95y31     80'h00_0060_00_0000_0C08_FFD3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1175_4 ( .OUT(na1175_2), .IN1(1'b0), .IN2(~na233_1), .IN3(~na1242_2), .IN4(na227_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x90y35     80'h00_0018_00_0000_0CEE_7500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1196_1 ( .OUT(na1196_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na232_1), .IN6(1'b0), .IN7(~na857_1), .IN8(~na227_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x88y31     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1198_4 ( .OUT(na1198_2), .IN1(1'b1), .IN2(~na261_2), .IN3(1'b1), .IN4(~na260_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y55     80'h00_0018_00_0040_0A55_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1200_1 ( .OUT(na1200_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na703_1), .IN4(1'b1), .IN5(~na670_2), .IN6(1'b0), .IN7(~na607_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x94y51     80'h00_0060_00_0000_0C08_FFB7
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1201_4 ( .OUT(na1201_2), .IN1(~na15_1), .IN2(~na1251_2), .IN3(na1200_1), .IN4(~na704_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y52     80'h00_0060_00_0000_0C08_FF58
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1203_4 ( .OUT(na1203_2), .IN1(na1219_2), .IN2(na7_2), .IN3(~na1201_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x73y128     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1204_4 ( .OUT(na1204_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na780_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1204_6 ( .RAM_O2(na1204_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1204_2), .COMP_OUT(1'b0) );
// C_///AND/      x75y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1205_4 ( .OUT(na1205_2), .IN1(na685_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1205_6 ( .RAM_O2(na1205_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1205_2), .COMP_OUT(1'b0) );
// C_///AND/      x77y128     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1206_4 ( .OUT(na1206_2), .IN1(1'b1), .IN2(na224_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1206_6 ( .RAM_O2(na1206_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1206_2), .COMP_OUT(1'b0) );
// C_///AND/      x115y1     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1207_4 ( .OUT(na1207_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na703_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1207_6 ( .RAM_O2(na1207_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1207_2), .COMP_OUT(1'b0) );
// C_///AND/      x113y1     80'h08_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1208_4 ( .OUT(na1208_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na704_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1208_6 ( .RAM_O2(na1208_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1208_2), .COMP_OUT(1'b0) );
// C_///AND/      x111y1     80'h08_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1209_4 ( .OUT(na1209_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na704_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1209_6 ( .RAM_O2(na1209_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1209_2), .COMP_OUT(1'b0) );
// C_///AND/      x109y1     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1210_4 ( .OUT(na1210_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na703_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1210_6 ( .RAM_O2(na1210_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1210_2), .COMP_OUT(1'b0) );
// C_///AND/      x107y1     80'h08_0060_00_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1211_4 ( .OUT(na1211_2), .IN1(~na707_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1211_6 ( .RAM_O2(na1211_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1211_2), .COMP_OUT(1'b0) );
// C_///AND/      x105y1     80'h08_0060_00_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1212_4 ( .OUT(na1212_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na708_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1212_6 ( .RAM_O2(na1212_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1212_2), .COMP_OUT(1'b0) );
// C_///AND/      x103y1     80'h08_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1213_4 ( .OUT(na1213_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na709_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1213_6 ( .RAM_O2(na1213_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1213_2), .COMP_OUT(1'b0) );
// C_///AND/      x101y1     80'h08_0060_00_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1214_4 ( .OUT(na1214_2), .IN1(1'b1), .IN2(~na710_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1214_6 ( .RAM_O2(na1214_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1214_2), .COMP_OUT(1'b0) );
// C_///AND/      x81y128     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1215_4 ( .OUT(na1215_2), .IN1(na788_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1215_6 ( .RAM_O2(na1215_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1215_2), .COMP_OUT(1'b0) );
// C_////Bridge      x89y44     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1216_5 ( .OUT(na1216_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1_1), .IN8(1'b0) );
// C_////Bridge      x94y53     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1217_5 ( .OUT(na1217_2), .IN1(na3_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1218_5 ( .OUT(na1218_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y51     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1219_5 ( .OUT(na1219_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na8_2), .IN8(1'b0) );
// C_////Bridge      x82y43     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1220_5 ( .OUT(na1220_2), .IN1(na10_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y58     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1221_5 ( .OUT(na1221_2), .IN1(na10_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y46     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1222_5 ( .OUT(na1222_2), .IN1(na10_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y61     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1223_5 ( .OUT(na1223_2), .IN1(na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y54     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1224_5 ( .OUT(na1224_2), .IN1(na10_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y43     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1225_5 ( .OUT(na1225_2), .IN1(1'b0), .IN2(1'b0), .IN3(na13_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y60     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1226_5 ( .OUT(na1226_2), .IN1(na18_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y37     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1227_5 ( .OUT(na1227_2), .IN1(1'b0), .IN2(na22_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y42     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1228_5 ( .OUT(na1228_2), .IN1(1'b0), .IN2(na22_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y49     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1229_5 ( .OUT(na1229_2), .IN1(1'b0), .IN2(na22_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x80y52     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1230_5 ( .OUT(na1230_2), .IN1(1'b0), .IN2(na22_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y62     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1231_5 ( .OUT(na1231_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na43_1) );
// C_////Bridge      x90y38     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1232_5 ( .OUT(na1232_2), .IN1(1'b0), .IN2(na46_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y54     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1233_5 ( .OUT(na1233_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na56_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y47     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1234_5 ( .OUT(na1234_2), .IN1(na93_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y49     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1235_5 ( .OUT(na1235_2), .IN1(na99_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y48     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1236_5 ( .OUT(na1236_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na107_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y57     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1237_5 ( .OUT(na1237_2), .IN1(na164_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y62     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1238_5 ( .OUT(na1238_2), .IN1(1'b0), .IN2(na170_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y61     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1239_5 ( .OUT(na1239_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na182_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y63     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1240_5 ( .OUT(na1240_2), .IN1(na189_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y65     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1241_5 ( .OUT(na1241_2), .IN1(na202_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y31     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1242_5 ( .OUT(na1242_2), .IN1(na232_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x94y29     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1243_5 ( .OUT(na1243_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na237_2) );
// C_////Bridge      x96y33     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1244_5 ( .OUT(na1244_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na241_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y29     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1245_5 ( .OUT(na1245_2), .IN1(1'b0), .IN2(na241_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y31     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1246_5 ( .OUT(na1246_2), .IN1(1'b0), .IN2(na245_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x85y31     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1247_5 ( .OUT(na1247_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na254_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y31     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1248_5 ( .OUT(na1248_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na260_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y29     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1249_5 ( .OUT(na1249_2), .IN1(na265_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x86y30     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1250_5 ( .OUT(na1250_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na265_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1251_5 ( .OUT(na1251_2), .IN1(1'b0), .IN2(1'b0), .IN3(na384_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y40     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1252_5 ( .OUT(na1252_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na428_1) );
// C_////Bridge      x93y40     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1253_5 ( .OUT(na1253_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na428_2) );
// C_////Bridge      x83y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1254_5 ( .OUT(na1254_2), .IN1(1'b0), .IN2(1'b0), .IN3(na447_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x82y48     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1255_5 ( .OUT(na1255_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na463_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x78y50     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1256_5 ( .OUT(na1256_2), .IN1(1'b0), .IN2(na465_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x87y30     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1257_5 ( .OUT(na1257_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na552_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y45     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1258_5 ( .OUT(na1258_2), .IN1(1'b0), .IN2(1'b0), .IN3(na568_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x83y47     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1259_5 ( .OUT(na1259_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na570_2) );
// C_////Bridge      x91y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1260_5 ( .OUT(na1260_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na592_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y57     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1261_5 ( .OUT(na1261_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na592_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y59     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1262_5 ( .OUT(na1262_2), .IN1(1'b0), .IN2(1'b0), .IN3(na612_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y65     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1263_5 ( .OUT(na1263_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na612_2), .IN8(1'b0) );
// C_////Bridge      x81y50     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1264_5 ( .OUT(na1264_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na631_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x81y48     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1265_5 ( .OUT(na1265_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na635_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y60     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1266_5 ( .OUT(na1266_2), .IN1(na657_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y58     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1267_5 ( .OUT(na1267_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na675_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y47     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1268_5 ( .OUT(na1268_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na703_1), .IN8(1'b0) );
// C_////Bridge      x95y48     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1269_5 ( .OUT(na1269_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na704_2) );
// C_////Bridge      x81y34     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1270_5 ( .OUT(na1270_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na920_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y50     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1271_5 ( .OUT(na1271_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na957_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y47     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1272_5 ( .OUT(na1272_2), .IN1(1'b0), .IN2(1'b0), .IN3(na962_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y48     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1273_5 ( .OUT(na1273_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na967_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y45     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1274_5 ( .OUT(na1274_2), .IN1(1'b0), .IN2(1'b0), .IN3(na972_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y46     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1275_5 ( .OUT(na1275_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na977_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y40     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1276_5 ( .OUT(na1276_2), .IN1(1'b0), .IN2(1'b0), .IN3(na980_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x77y43     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1277_5 ( .OUT(na1277_2), .IN1(1'b0), .IN2(1'b0), .IN3(na983_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y44     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1278_5 ( .OUT(na1278_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na989_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x79y43     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1279_5 ( .OUT(na1279_2), .IN1(1'b0), .IN2(1'b0), .IN3(na992_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y48     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1280_5 ( .OUT(na1280_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1030_1) );
// C_////Bridge      x90y53     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1281_5 ( .OUT(na1281_2), .IN1(1'b0), .IN2(na1152_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y63     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1282_5 ( .OUT(na1282_2), .IN1(1'b0), .IN2(na1165_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
endmodule
