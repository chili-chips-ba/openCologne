//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 July 2024)
//  Compile Time: 1970-01-01 00:59:59
//  Program Run:  2024-07-21 11:15:13
//  Program Call: p_r +sp -i /home/user/openCologne/1.Blinky--ILA-Test/net/ila_top_synth24-07-21_11-14-53.v -o /home/user/openCologne/1.Blinky--ILA-Test/p_r_out/ila_top_24-07-21_11-14-53 -sp -cCP +uCIO -ccf /home/user/openCologne/1.Blinky--ILA-Test/src/ILA_top.ccf 
//  File Type:    Verilog

// Gatecount:    263
module ila_top_24-07-21_11-14-53 (clk , i_mosi_ILA , i_sclk_ILA , i_ss_ILA ,
       led , o_miso_ILA 
       ) ;

input  clk;
input  i_mosi_ILA;
input  i_sclk_ILA;
input  i_ss_ILA;

output led;
output o_miso_ILA;



wire clk;
wire led;
wire na1_1;
wire na1_1_i;
wire na1_2;
wire na1_2_i;
wire na2_1;
wire na2_1_i;
wire na3_1;
wire na4_1;
wire na4_1_i;
wire na4_2;
wire na4_2_i;
wire na5_1;
wire na5_1_i;
wire na6_2;
wire na6_2_i;
wire na7_1;
wire na8_1;
wire na8_1_i;
wire na8_2;
wire na8_2_i;
wire na9_1;
wire na9_1_i;
wire na9_2;
wire na9_2_i;
wire na10_1;
wire na10_1_i;
wire na13_1;
wire na13_1_i;
wire na13_2;
wire na13_2_i;
wire na15_1;
wire na15_1_i;
wire na15_2;
wire na15_2_i;
wire na16_1;
wire na16_1_i;
wire na16_2;
wire na16_2_i;
wire na17_1;
wire na17_1_i;
wire na17_2;
wire na17_2_i;
wire na19_1;
wire na19_1_i;
wire na20_1;
wire na20_1_i;
wire na21_2;
wire na21_2_i;
wire na22_2;
wire na24_1;
wire na24_1_i;
wire na24_2;
wire na24_2_i;
wire na25_1;
wire na25_1_i;
wire na25_2;
wire na25_2_i;
wire na26_1;
wire na26_1_i;
wire na26_2;
wire na26_2_i;
wire na27_1;
wire na27_1_i;
wire na27_2;
wire na27_2_i;
wire na31_1;
wire na31_1_i;
wire na31_2;
wire na31_2_i;
wire na32_1;
wire na32_1_i;
wire na33_1;
wire na33_1_i;
wire na34_2;
wire na34_2_i;
wire na35_1;
wire na35_1_i;
wire na36_1;
wire na36_1_i;
wire na36_2;
wire na36_2_i;
wire na37_1;
wire na37_1_i;
wire na37_2;
wire na37_2_i;
wire na38_1;
wire na38_1_i;
wire na40_1;
wire na40_1_i;
wire na40_2;
wire na40_2_i;
wire na42_2;
wire na42_2_i;
wire na43_1;
wire na43_1_i;
wire na43_2;
wire na43_2_i;
wire na44_1;
wire na44_1_i;
wire na45_1;
wire na45_1_i;
wire na47_1;
wire na47_1_i;
wire na47_2;
wire na47_2_i;
wire na49_1;
wire na49_1_i;
wire na49_2;
wire na49_2_i;
wire na51_1;
wire na51_1_i;
wire na51_2;
wire na51_2_i;
wire na53_2;
wire na53_2_i;
wire na54_2;
wire na55_1;
wire na55_1_i;
wire na55_2;
wire na55_2_i;
wire na56_1;
wire na56_1_i;
wire na56_2;
wire na56_2_i;
wire na58_1;
wire na58_1_i;
wire na59_1;
wire na60_2;
wire na60_2_i;
wire na61_1;
wire na61_1_i;
wire na62_1;
wire na62_1_i;
wire na62_2;
wire na62_2_i;
wire na63_1;
wire na63_1_i;
wire na63_2;
wire na63_2_i;
wire na67_1;
wire na67_1_i;
wire na67_2;
wire na67_2_i;
wire na70_1;
wire na70_1_i;
wire na73_1;
wire na73_1_i;
wire na73_2;
wire na73_2_i;
wire na75_1;
wire na75_1_i;
wire na76_1;
wire na76_1_i;
wire na78_1;
wire na78_1_i;
wire na78_2;
wire na78_2_i;
wire na79_1;
wire na79_1_i;
wire na79_2;
wire na79_2_i;
wire na83_1;
wire na83_1_i;
wire na87_1;
wire na87_1_i;
wire na88_1;
wire na88_1_i;
wire na89_1;
wire na89_1_i;
wire na90_1;
wire na90_1_i;
wire na91_1;
wire na91_1_i;
wire na92_1;
wire na92_1_i;
wire na93_1;
wire na93_1_i;
wire na94_1;
wire na94_1_i;
wire na95_1;
wire na95_1_i;
wire na97_1;
wire na97_1_i;
wire na100_1;
wire na100_1_i;
wire na100_2;
wire na100_2_i;
wire na101_1;
wire na101_1_i;
wire na101_2;
wire na101_2_i;
wire na104_1;
wire na104_1_i;
wire na106_2;
wire na106_2_i;
wire na107_1;
wire na107_1_i;
wire na108_1;
wire na108_1_i;
wire na108_2;
wire na108_2_i;
wire na109_1;
wire na109_1_i;
wire na110_1;
wire na110_1_i;
wire na111_1;
wire na111_1_i;
wire na111_2;
wire na111_2_i;
wire na112_2;
wire na112_2_i;
wire na113_1;
wire na113_1_i;
wire na115_2;
wire na115_2_i;
wire na116_2;
wire na120_1;
wire na121_1;
wire na121_1_i;
wire na122_1;
wire na123_1;
wire na123_1_i;
wire na126_1;
wire na126_2;
wire na126_4;
wire na128_1;
wire na128_2;
wire na128_4;
wire na130_1;
wire na130_2;
wire na130_4;
wire na132_1;
wire na132_2;
wire na132_4;
wire na134_1;
wire na134_2;
wire na134_4;
wire na135_1;
wire na135_2;
wire na135_4;
wire na137_1;
wire na137_2;
wire na137_4;
wire na139_1;
wire na139_2;
wire na142_1;
wire na142_2;
wire na142_4;
wire na144_1;
wire na144_2;
wire na144_4;
wire na146_1;
wire na146_2;
wire na146_4;
wire na148_1;
wire na148_2;
wire na148_4;
wire na149_1;
wire na149_4;
wire na150_1;
wire na150_2;
wire na150_4;
wire na152_1;
wire na152_2;
wire na152_4;
wire na154_1;
wire na154_2;
wire na154_4;
wire na156_1;
wire na156_2;
wire na158_1;
wire na158_4;
wire na159_1;
wire na159_2;
wire na159_4;
wire na161_1;
wire na161_2;
wire na161_4;
wire na163_1;
wire na163_2;
wire na163_4;
wire na165_1;
wire na165_2;
wire na167_1;
wire na167_4;
wire na168_1;
wire na168_2;
wire na168_4;
wire na170_1;
wire na170_2;
wire na170_4;
wire na172_1;
wire na172_2;
wire na172_4;
wire na174_1;
wire na174_2;
wire na176_1;
wire na176_4;
wire na177_1;
wire na177_2;
wire na177_4;
wire na179_1;
wire na179_2;
wire na179_4;
wire na181_1;
wire na181_2;
wire na181_4;
wire na183_1;
wire na183_2;
wire na187_1;
wire na187_2;
wire na204_1;
wire na204_1_i;
wire na205_2;
wire na205_2_i;
wire na255_1;
wire na255_1_i;
wire na265_2;
wire na265_2_i;
wire na298_1;
wire na299_1;
wire na300_1;
wire na301_1;
wire na304_3;
wire na304_4;
wire na304_5;
wire na304_6;
wire na305_3;
wire na305_4;
wire na305_5;
wire na305_6;
wire na307_1;
wire na308_1;
wire na308_2;
wire na309_1;
wire na310_1;
wire na311_1;
wire na312_2;
wire na313_1;
wire na313_9;
wire na314_2;
wire na315_1;
wire na316_1;
wire na317_1;
wire na318_1;
wire na319_2;
wire na320_1;
wire na321_1;
wire na322_1;
wire na323_1;
wire na324_1;
wire na325_1;
wire na326_1;
wire na326_9;
wire na327_1;
wire na328_1;
wire na329_1;
wire na330_1;
wire na331_1;
wire na332_1;
wire na333_2;
wire na334_2;
wire na335_1;
wire na336_1;
wire na336_9;
wire na337_2;
wire na338_2;
wire na339_1;
wire na339_4;
wire na340_1;
wire na340_9;
wire na341_2;
wire na342_1;
wire na342_9;
wire na343_1;
wire na344_2;
wire na345_1;
wire na345_9;
wire na346_2;
wire na347_1;
wire na348_1;
wire na349_1;
wire na350_1;
wire na351_1;
wire na351_9;
wire na352_1;
wire na353_2;
wire na354_1;
wire na355_1;
wire na356_1;
wire na357_1;
wire na358_1;
wire na359_1;
wire na359_9;
wire na360_2;
wire na361_1;
wire na362_1;
wire na363_1;
wire na364_1;
wire na364_9;
wire na365_1;
wire na366_2;
wire na367_1;
wire na367_9;
wire na368_2;
wire na369_2;
wire na370_2;
wire na371_2;
wire na372_1;
wire na372_9;
wire na373_2;
wire na374_1;
wire na374_9;
wire na375_2;
wire na376_1;
wire na376_9;
wire na377_2;
wire na378_1;
wire na378_9;
wire na379_2;
wire na380_1;
wire na380_9;
wire na381_2;
wire na382_1;
wire na382_9;
wire na383_2;
wire na384_1;
wire na384_9;
wire na385_2;
wire na386_1;
wire na386_9;
wire na387_2;
wire na388_1;
wire na388_9;
wire na389_2;
wire na390_1;
wire na390_9;
wire na391_2;
wire na392_1;
wire na392_9;
wire na393_2;
wire na394_1;
wire na394_9;
wire na395_2;
wire na396_1;
wire na396_9;
wire na397_2;
wire na398_1;
wire na398_9;
wire na399_2;
wire na400_1;
wire na400_9;
wire na401_2;
wire na402_1;
wire na402_9;
wire na403_2;
wire na404_1;
wire na404_9;
wire na405_2;
wire na406_1;
wire na406_9;
wire na407_2;
wire na408_1;
wire na408_9;
wire na409_2;
wire na410_1;
wire na410_9;
wire na411_2;
wire na412_1;
wire na412_9;
wire na413_2;
wire na414_1;
wire na414_9;
wire na415_2;
wire na416_1;
wire na416_9;
wire na417_2;
wire na418_1;
wire na418_9;
wire na419_2;
wire na420_1;
wire na421_2;
wire na422_2;
wire na423_2;
wire na424_2;
wire na425_2;
wire na426_2;
wire na427_2;
wire na428_2;
wire na429_2;
wire na430_2;
wire na431_2;
wire na432_2;
wire na433_2;
wire na434_2;
wire na435_2;
wire na436_2;
wire na437_2;
wire na438_2;
wire na439_2;
wire na440_2;
wire na441_2;
wire na442_2;
wire na443_2;
wire na444_2;
wire na445_2;
wire na446_2;
wire i_ss_ILA;
wire na314_10;
wire na319_10;
wire na333_10;
wire na338_10;
wire na341_10;
wire na344_10;
wire na346_10;
wire na353_10;
wire na360_10;
wire na366_10;
wire na369_10;
wire na370_10;
wire na371_10;
wire na373_10;
wire na375_10;
wire na377_10;
wire na379_10;
wire na381_10;
wire na383_10;
wire na385_10;
wire na387_10;
wire na389_10;
wire na391_10;
wire na393_10;
wire na395_10;
wire na397_10;
wire na399_10;
wire na401_10;
wire na403_10;
wire na405_10;
wire na407_10;
wire na409_10;
wire na411_10;
wire na413_10;
wire na415_10;
wire na417_10;
wire na419_10;
wire na306_120;
wire i_mosi_ILA;
wire i_sclk_ILA;
wire o_miso_ILA;

// C_ICOMP/D//AND/D      x12y35     80'h00_FE00_80_0000_0C88_6A82
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1_1 ( .OUT(na1_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na109_1), .IN6(1'b0), .IN7(na1_2), .IN8(~na421_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1_2 ( .OUT(na1_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1_4 ( .OUT(na1_2_i), .IN1(na109_1), .IN2(~na433_2), .IN3(na19_1), .IN4(na443_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1_5 ( .OUT(na1_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1_2_i) );
// C_MX4b/D///      x17y38     80'h00_FD00_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a2_1 ( .OUT(na2_1_i), .IN1(~na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(na301_1), .IN5(na9_2), .IN6(na2_1), .IN7(1'b0), .IN8(1'b0),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2_2 ( .OUT(na2_1), .CLK(~na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2_1_i) );
// C_AND////      x17y35     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3_1 ( .OUT(na3_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na435_2), .IN7(1'b1), .IN8(na73_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x8y45     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4_1 ( .OUT(na4_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na126_2), .IN6(na312_2), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a4_2 ( .OUT(na4_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4_4 ( .OUT(na4_2_i), .IN1(na126_1), .IN2(na312_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a4_5 ( .OUT(na4_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na4_2_i) );
// C_AND/D///      x16y38     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a5_1 ( .OUT(na5_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(1'b1), .IN7(na309_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a5_2 ( .OUT(na5_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na5_1_i) );
// C_///AND/D      x17y36     80'h00_FD00_80_0000_0C08_FF1A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6_4 ( .OUT(na6_2_i), .IN1(na3_1), .IN2(1'b1), .IN3(~na7_1), .IN4(~na301_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6_5 ( .OUT(na6_2), .CLK(~na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6_2_i) );
// C_MX2b////      x16y37     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a7_1 ( .OUT(na7_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na55_2), .IN5(~na9_1), .IN6(1'b0), .IN7(~na310_1), .IN8(1'b0),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x11y42     80'h00_FE00_80_0000_0C88_ACA2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na8_2), .IN7(na75_1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a8_2 ( .OUT(na8_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na8_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a8_4 ( .OUT(na8_2_i), .IN1(na83_1), .IN2(~na15_2), .IN3(na75_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a8_5 ( .OUT(na8_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na8_2_i) );
// C_AND/D//AND/D      x15y37     80'h00_FE00_80_0000_0C88_3C3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9_1 ( .OUT(na9_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na299_1), .IN7(1'b1), .IN8(~na301_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a9_2 ( .OUT(na9_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na9_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9_4 ( .OUT(na9_2_i), .IN1(na9_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na301_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a9_5 ( .OUT(na9_2), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na9_2_i) );
// C_AND/D///      x17y40     80'h00_FE00_00_0000_0888_A12C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a10_1 ( .OUT(na10_1_i), .IN1(1'b1), .IN2(na34_2), .IN3(na61_1), .IN4(~na33_1), .IN5(~na44_1), .IN6(~na2_1), .IN7(na35_1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a10_2 ( .OUT(na10_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na10_1_i) );
// C_AND/D//AND/D      x8y46     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na139_2), .IN6(na312_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a13_2 ( .OUT(na13_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na13_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a13_4 ( .OUT(na13_2_i), .IN1(na139_1), .IN2(na312_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a13_5 ( .OUT(na13_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na13_2_i) );
// C_AND/D//AND/D      x11y44     80'h00_FE00_80_0000_0C88_A4FC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a15_1 ( .OUT(na15_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na83_1), .IN6(na15_2), .IN7(na75_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a15_2 ( .OUT(na15_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na15_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a15_4 ( .OUT(na15_2_i), .IN1(1'b1), .IN2(na101_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a15_5 ( .OUT(na15_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na15_2_i) );
// C_AND/D//AND/D      x22y33     80'h00_FE00_80_0000_0C88_3A2F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a16_1 ( .OUT(na16_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na9_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na301_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a16_2 ( .OUT(na16_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na16_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a16_4 ( .OUT(na16_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na16_1), .IN4(~na301_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a16_5 ( .OUT(na16_2), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na16_2_i) );
// C_AND/D//AND/D      x16y34     80'h00_FE00_80_0000_0C88_2AAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a17_1 ( .OUT(na17_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(1'b1), .IN7(na265_2), .IN8(~na17_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a17_2 ( .OUT(na17_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na17_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a17_4 ( .OUT(na17_2_i), .IN1(na109_1), .IN2(1'b1), .IN3(na320_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a17_5 ( .OUT(na17_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na17_2_i) );
// C_ORAND/D///      x14y33     80'h00_FE00_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a19_1 ( .OUT(na19_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(1'b0), .IN7(na19_1), .IN8(na17_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a19_2 ( .OUT(na19_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na19_1_i) );
// C_ORAND/D///      x15y40     80'h00_FE00_00_0000_0888_FE5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a20_1 ( .OUT(na20_1_i), .IN1(1'b0), .IN2(na312_2), .IN3(~na97_1), .IN4(1'b0), .IN5(na204_1), .IN6(na20_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a20_2 ( .OUT(na20_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na20_1_i) );
// C_///ICOMP/D      x16y45     80'h00_FE00_80_0000_0C08_FF6C
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a21_4 ( .OUT(na21_2_i), .IN1(1'b0), .IN2(~na20_1), .IN3(na21_2), .IN4(~na22_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a21_5 ( .OUT(na21_2), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na21_2_i) );
// C_///AND/      x18y40     80'h00_0060_00_0000_0C08_FFC8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a22_4 ( .OUT(na22_2), .IN1(na44_1), .IN2(na32_1), .IN3(1'b1), .IN4(na429_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//ORAND/D      x15y39     80'h00_FE00_80_0000_0C88_AAEC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a24_1 ( .OUT(na24_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na24_2), .IN6(1'b1), .IN7(na420_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a24_2 ( .OUT(na24_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na24_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a24_4 ( .OUT(na24_2_i), .IN1(1'b0), .IN2(na20_1), .IN3(na334_2), .IN4(na428_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a24_5 ( .OUT(na24_2), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na24_2_i) );
// C_AND/D//AND/D      x15y32     80'h00_FE00_80_0000_0C88_AACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a25_1 ( .OUT(na25_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(1'b1), .IN7(na315_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a25_2 ( .OUT(na25_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na25_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a25_4 ( .OUT(na25_2_i), .IN1(na109_1), .IN2(1'b1), .IN3(1'b1), .IN4(na316_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a25_5 ( .OUT(na25_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na25_2_i) );
// C_AND/D//AND/D      x8y43     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a26_1 ( .OUT(na26_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na132_2), .IN7(na444_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a26_2 ( .OUT(na26_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na26_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a26_4 ( .OUT(na26_2_i), .IN1(1'b1), .IN2(na132_1), .IN3(na444_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a26_5 ( .OUT(na26_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na26_2_i) );
// C_AND/D//AND/D      x9y46     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na137_2), .IN7(na444_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a27_2 ( .OUT(na27_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na27_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a27_4 ( .OUT(na27_2_i), .IN1(1'b1), .IN2(na137_1), .IN3(na444_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a27_5 ( .OUT(na27_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na27_2_i) );
// C_AND/D//AND/D      x10y46     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a31_1 ( .OUT(na31_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na134_2), .IN6(na312_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a31_2 ( .OUT(na31_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na31_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a31_4 ( .OUT(na31_2_i), .IN1(na134_1), .IN2(na312_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a31_5 ( .OUT(na31_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na31_2_i) );
// C_MX4a/D///      x17y42     80'h00_FE00_00_0040_0C0A_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a32_1 ( .OUT(na32_1_i), .IN1(1'b0), .IN2(na32_1), .IN3(1'b0), .IN4(na317_1), .IN5(1'b1), .IN6(na20_1), .IN7(1'b1), .IN8(na430_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a32_2 ( .OUT(na32_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na32_1_i) );
// C_MX4b/D///      x16y42     80'h00_FD00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_1 ( .OUT(na33_1_i), .IN1(~na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na301_1), .IN5(1'b0), .IN6(1'b0), .IN7(na16_1), .IN8(na33_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a33_2 ( .OUT(na33_1), .CLK(~na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na33_1_i) );
// C_///AND/D      x21y36     80'h00_FD00_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a34_4 ( .OUT(na34_2_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na301_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a34_5 ( .OUT(na34_2), .CLK(~na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na34_2_i) );
// C_MX4b/D///      x18y41     80'h00_FD00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a35_1 ( .OUT(na35_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na301_1), .IN5(1'b0), .IN6(1'b0), .IN7(na35_1), .IN8(na425_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a35_2 ( .OUT(na35_1), .CLK(~na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na35_1_i) );
// C_AND/D//AND/D      x8y42     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na130_2), .IN6(na312_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a36_2 ( .OUT(na36_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na36_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a36_4 ( .OUT(na36_2_i), .IN1(na130_1), .IN2(na312_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a36_5 ( .OUT(na36_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na36_2_i) );
// C_AND/D//AND/D      x7y45     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a37_1 ( .OUT(na37_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na146_2), .IN6(na312_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a37_2 ( .OUT(na37_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na37_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a37_4 ( .OUT(na37_2_i), .IN1(na146_1), .IN2(na312_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a37_5 ( .OUT(na37_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na37_2_i) );
// C_AND/D///      x14y36     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a38_1 ( .OUT(na38_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na318_1), .IN6(1'b1), .IN7(1'b1), .IN8(na442_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a38_2 ( .OUT(na38_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na38_1_i) );
// C_AND/D//AND/D      x7y43     80'h00_FE00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a40_1 ( .OUT(na40_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na142_2), .IN6(na312_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a40_2 ( .OUT(na40_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na40_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a40_4 ( .OUT(na40_2_i), .IN1(na142_1), .IN2(na312_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a40_5 ( .OUT(na40_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na40_2_i) );
// C_///AND/D      x10y43     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a42_4 ( .OUT(na42_2_i), .IN1(na445_2), .IN2(na135_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a42_5 ( .OUT(na42_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na42_2_i) );
// C_AND/D//AND/D      x14y35     80'h00_FE00_80_0000_0C88_4ACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a43_1 ( .OUT(na43_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(1'b1), .IN7(~na43_2), .IN8(na255_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a43_2 ( .OUT(na43_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na43_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a43_4 ( .OUT(na43_2_i), .IN1(na109_1), .IN2(1'b1), .IN3(1'b1), .IN4(na355_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a43_5 ( .OUT(na43_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na43_2_i) );
// C_ORAND/D///      x15y35     80'h00_FE00_00_0000_0888_FEA5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a44_1 ( .OUT(na44_1_i), .IN1(~na109_1), .IN2(1'b0), .IN3(na426_2), .IN4(1'b0), .IN5(na44_1), .IN6(na10_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a44_2 ( .OUT(na44_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na44_1_i) );
// C_AND/D///      x21y39     80'h00_FE00_00_0000_0888_A344
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1_i), .IN1(~na44_1), .IN2(na34_2), .IN3(~na61_1), .IN4(na33_1), .IN5(1'b1), .IN6(~na2_1), .IN7(na35_1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a45_2 ( .OUT(na45_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na45_1_i) );
// C_AND/D//AND/D      x11y46     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a47_1 ( .OUT(na47_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na148_2), .IN7(na444_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a47_2 ( .OUT(na47_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na47_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a47_4 ( .OUT(na47_2_i), .IN1(1'b1), .IN2(na148_1), .IN3(na444_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a47_5 ( .OUT(na47_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na47_2_i) );
// C_AND/D//AND/D      x15y34     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a49_1 ( .OUT(na49_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(1'b1), .IN7(na321_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a49_2 ( .OUT(na49_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na49_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a49_4 ( .OUT(na49_2_i), .IN1(na109_1), .IN2(1'b1), .IN3(na322_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a49_5 ( .OUT(na49_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na49_2_i) );
// C_AND/D//AND/D      x15y31     80'h00_FE00_80_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a51_1 ( .OUT(na51_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(1'b1), .IN7(na323_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a51_2 ( .OUT(na51_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na51_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a51_4 ( .OUT(na51_2_i), .IN1(na109_1), .IN2(na324_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a51_5 ( .OUT(na51_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na51_2_i) );
// C_///AND/D      x14y41     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a53_4 ( .OUT(na53_2_i), .IN1(1'b1), .IN2(na20_1), .IN3(1'b1), .IN4(na325_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a53_5 ( .OUT(na53_2), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na53_2_i) );
// C_///AND/      x15y42     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a54_4 ( .OUT(na54_2), .IN1(na44_1), .IN2(na32_1), .IN3(na21_2), .IN4(na429_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP/D//ORAND/D      x16y32     80'h00_FE00_80_0000_0C88_9AEA
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na109_1), .IN6(1'b0), .IN7(~na432_2), .IN8(~na55_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a55_2 ( .OUT(na55_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na55_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a55_4 ( .OUT(na55_2_i), .IN1(na109_1), .IN2(1'b0), .IN3(na43_1), .IN4(na55_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a55_5 ( .OUT(na55_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na55_2_i) );
// C_AND/D//AND/D      x21y35     80'h00_FE00_80_0000_0C88_F8AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a56_1 ( .OUT(na56_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(na327_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a56_2 ( .OUT(na56_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na56_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a56_4 ( .OUT(na56_2_i), .IN1(na109_1), .IN2(1'b1), .IN3(na328_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a56_5 ( .OUT(na56_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na56_2_i) );
// C_AND/D///      x14y41     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a58_1 ( .OUT(na58_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na329_1), .IN6(na20_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a58_2 ( .OUT(na58_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na58_1_i) );
// C_AND////      x15y41     80'h00_0018_00_0000_0C88_82FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a59_1 ( .OUT(na59_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na44_1), .IN6(~na32_1), .IN7(na21_2), .IN8(na429_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x16y44     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a60_4 ( .OUT(na60_2_i), .IN1(1'b1), .IN2(na20_1), .IN3(na330_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a60_5 ( .OUT(na60_2), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na60_2_i) );
// C_MX4b/D///      x16y41     80'h00_FD00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a61_1 ( .OUT(na61_1_i), .IN1(na3_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na301_1), .IN5(1'b0), .IN6(1'b0), .IN7(na61_1), .IN8(na423_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a61_2 ( .OUT(na61_1), .CLK(~na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na61_1_i) );
// C_AND/D//AND/D      x7y46     80'h00_FE00_80_0000_0C88_ACA3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a62_1 ( .OUT(na62_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na135_2), .IN7(na444_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a62_2 ( .OUT(na62_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na62_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a62_4 ( .OUT(na62_2_i), .IN1(1'b1), .IN2(~na62_2), .IN3(na444_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a62_5 ( .OUT(na62_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na62_2_i) );
// C_AND/D//AND/D      x11y45     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a63_1 ( .OUT(na63_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na144_2), .IN7(na444_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a63_2 ( .OUT(na63_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na63_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a63_4 ( .OUT(na63_2_i), .IN1(1'b1), .IN2(na144_1), .IN3(na444_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a63_5 ( .OUT(na63_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na63_2_i) );
// C_AND/D//AND/D      x20y33     80'h00_FE00_80_0000_0C88_AAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_1 ( .OUT(na67_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(1'b1), .IN7(na331_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a67_2 ( .OUT(na67_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na67_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a67_4 ( .OUT(na67_2_i), .IN1(na109_1), .IN2(na332_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a67_5 ( .OUT(na67_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na67_2_i) );
// C_ORAND/D///      x14y32     80'h00_FD00_00_0000_0888_3F3E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a70_1 ( .OUT(na70_1_i), .IN1(na3_1), .IN2(na6_2), .IN3(1'b0), .IN4(~na335_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0), .IN8(~na301_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a70_2 ( .OUT(na70_1), .CLK(~na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na70_1_i) );
// C_AND*/D//ICOMP*/D      x22y38     80'h00_FE00_80_0000_0387_C339
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a73_1 ( .OUT(na73_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na301_1), .IN7(1'b1), .IN8(na73_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a73_2 ( .OUT(na73_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na73_1_i) );
C_ICOMP    #(.CPE_CFG (9'b1_1000_0000)) 
           _a73_4 ( .OUT(na73_2_i), .IN1(~na436_2), .IN2(~na435_2), .IN3(1'b0), .IN4(na301_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a73_5 ( .OUT(na73_2), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na73_2_i) );
// C_ORAND/D///      x14y45     80'h00_FE00_00_0000_0888_EF5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1_i), .IN1(1'b0), .IN2(na312_2), .IN3(~na97_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na75_1), .IN8(na205_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a75_2 ( .OUT(na75_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na75_1_i) );
// C_ORAND/D///      x17y27     80'h00_FD00_00_0000_0888_3F3E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a76_1 ( .OUT(na76_1_i), .IN1(na3_1), .IN2(na121_1), .IN3(1'b0), .IN4(~na343_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0), .IN8(~na301_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a76_2 ( .OUT(na76_1), .CLK(~na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na76_1_i) );
// C_AND/D//AND/D      x14y37     80'h00_FE00_80_0000_0C88_CAF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(1'b1), .IN7(1'b1), .IN8(na347_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a78_2 ( .OUT(na78_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a78_4 ( .OUT(na78_2_i), .IN1(na109_1), .IN2(na311_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a78_5 ( .OUT(na78_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_2_i) );
// C_AND/D//AND/D      x21y31     80'h00_FE00_80_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a79_1 ( .OUT(na79_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na348_1), .IN6(1'b1), .IN7(1'b1), .IN8(na442_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a79_2 ( .OUT(na79_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na79_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a79_4 ( .OUT(na79_2_i), .IN1(na109_1), .IN2(1'b1), .IN3(1'b1), .IN4(na352_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a79_5 ( .OUT(na79_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na79_2_i) );
// C_MX2b/D///      x15y45     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a83_1 ( .OUT(na83_1_i), .IN1(1'b1), .IN2(na438_2), .IN3(1'b0), .IN4(1'b0), .IN5(na439_2), .IN6(na15_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a83_2 ( .OUT(na83_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na83_1_i) );
// C_MX2b/D///      x20y34     80'h00_FA00_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a87_1 ( .OUT(na87_1_i), .IN1(1'b1), .IN2(na34_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na111_2), .IN8(~na87_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a87_2 ( .OUT(na87_1), .CLK(na300_1), .EN(na116_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na87_1_i) );
// C_MX2b/D///      x19y36     80'h00_FA00_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a88_1 ( .OUT(na88_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_2), .IN5(1'b0), .IN6(na150_1), .IN7(1'b0), .IN8(na159_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a88_2 ( .OUT(na88_1), .CLK(na300_1), .EN(na116_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na88_1_i) );
// C_MX2b/D///      x20y35     80'h00_FA00_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_2), .IN5(1'b0), .IN6(na150_2), .IN7(1'b0), .IN8(na159_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a89_2 ( .OUT(na89_1), .CLK(na300_1), .EN(na116_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_1_i) );
// C_MX2b/D///      x20y36     80'h00_FA00_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_2), .IN5(na152_1), .IN6(1'b0), .IN7(na161_1), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a90_2 ( .OUT(na90_1), .CLK(na300_1), .EN(na116_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na90_1_i) );
// C_MX2b/D///      x17y37     80'h00_FA00_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a91_1 ( .OUT(na91_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_2), .IN5(na152_2), .IN6(1'b0), .IN7(na161_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a91_2 ( .OUT(na91_1), .CLK(na300_1), .EN(na116_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na91_1_i) );
// C_MX2b/D///      x16y39     80'h00_FA00_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a92_1 ( .OUT(na92_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_2), .IN5(1'b0), .IN6(na154_1), .IN7(1'b0), .IN8(na163_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a92_2 ( .OUT(na92_1), .CLK(na300_1), .EN(na116_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na92_1_i) );
// C_MX2b/D///      x17y39     80'h00_FA00_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_1 ( .OUT(na93_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na429_2), .IN5(1'b0), .IN6(na154_2), .IN7(1'b0), .IN8(na163_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a93_2 ( .OUT(na93_1), .CLK(na300_1), .EN(na116_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na93_1_i) );
// C_MX2b/D///      x18y39     80'h00_FA00_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a94_1 ( .OUT(na94_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_2), .IN5(na156_1), .IN6(1'b0), .IN7(na165_1), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a94_2 ( .OUT(na94_1), .CLK(na300_1), .EN(na116_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na94_1_i) );
// C_MX2b/D///      x20y40     80'h00_FA00_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a95_1 ( .OUT(na95_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na429_2), .IN5(na156_2), .IN6(1'b0), .IN7(na165_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a95_2 ( .OUT(na95_1), .CLK(na300_1), .EN(na116_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na95_1_i) );
// C_AND/D///      x18y43     80'h00_FE00_00_0000_0888_4C54
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a97_1 ( .OUT(na97_1_i), .IN1(~na44_1), .IN2(na34_2), .IN3(~na61_1), .IN4(1'b1), .IN5(1'b1), .IN6(na2_1), .IN7(~na35_1),
                    .IN8(na33_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a97_2 ( .OUT(na97_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na97_1_i) );
// C_AND/D//AND/D      x13y46     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a100_1 ( .OUT(na100_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na128_2), .IN7(na444_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a100_2 ( .OUT(na100_1), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na100_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a100_4 ( .OUT(na100_2_i), .IN1(1'b1), .IN2(na128_1), .IN3(na444_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a100_5 ( .OUT(na100_2), .CLK(na187_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na100_2_i) );
// C_AND/D//AND/D      x15y46     80'h00_FE00_80_0000_0C88_14AA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a101_1 ( .OUT(na101_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na104_1), .IN6(na101_2), .IN7(~na58_1), .IN8(~na60_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a101_2 ( .OUT(na101_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na101_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a101_4 ( .OUT(na101_2_i), .IN1(na298_1), .IN2(1'b1), .IN3(na75_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a101_5 ( .OUT(na101_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na101_2_i) );
// C_AND/D///      x15y43     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a104_1 ( .OUT(na104_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na20_1), .IN7(1'b1), .IN8(na354_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a104_2 ( .OUT(na104_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na104_1_i) );
// C_///AND/D      x14y33     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a106_4 ( .OUT(na106_2_i), .IN1(na109_1), .IN2(na356_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a106_5 ( .OUT(na106_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na106_2_i) );
// C_AND/D///      x18y42     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a107_1 ( .OUT(na107_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na20_1), .IN7(na357_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a107_2 ( .OUT(na107_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na107_1_i) );
// C_AND/D//AND/D      x14y34     80'h00_FE00_80_0000_0C88_F8CA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a108_1 ( .OUT(na108_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(na358_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a108_2 ( .OUT(na108_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na108_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a108_4 ( .OUT(na108_2_i), .IN1(na109_1), .IN2(1'b1), .IN3(1'b1), .IN4(na350_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a108_5 ( .OUT(na108_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na108_2_i) );
// C_ORAND/D///      x13y31     80'h00_FE00_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a109_1 ( .OUT(na109_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(na54_2), .IN7(1'b0), .IN8(na427_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a109_2 ( .OUT(na109_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na109_1_i) );
// C_ORAND/D///      x21y38     80'h00_FE00_00_0000_0888_FE3C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a110_1 ( .OUT(na110_1_i), .IN1(1'b0), .IN2(na20_1), .IN3(1'b0), .IN4(~na428_2), .IN5(na45_1), .IN6(na110_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a110_2 ( .OUT(na110_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na110_1_i) );
// C_AND/D//AND/D      x20y31     80'h00_FE00_80_0000_0C88_AAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a111_1 ( .OUT(na111_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na109_1), .IN6(1'b1), .IN7(na361_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a111_2 ( .OUT(na111_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na111_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a111_4 ( .OUT(na111_2_i), .IN1(na109_1), .IN2(1'b1), .IN3(na349_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a111_5 ( .OUT(na111_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na111_2_i) );
// C_///OR/D      x10y34     80'h00_FE00_80_0000_0C0E_FFC5
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a112_4 ( .OUT(na112_2_i), .IN1(~na109_1), .IN2(1'b0), .IN3(1'b0), .IN4(na362_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a112_5 ( .OUT(na112_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na112_2_i) );
// C_AND/D///      x12y44     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a113_1 ( .OUT(na113_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na15_1), .IN7(na75_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a113_2 ( .OUT(na113_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na113_1_i) );
// C_///AND/D      x23y34     80'h00_FE00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a115_4 ( .OUT(na115_2_i), .IN1(na109_1), .IN2(1'b1), .IN3(1'b1), .IN4(na363_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a115_5 ( .OUT(na115_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na115_2_i) );
// C_///OR/      x20y37     80'h00_0060_00_0000_0C0E_FFAC
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a116_4 ( .OUT(na116_2), .IN1(1'b0), .IN2(na34_2), .IN3(na337_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x13y38     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a120_1 ( .OUT(na120_1), .IN1(1'b1), .IN2(na433_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na16_1), .IN8(~na365_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x19y32     80'h00_FD00_00_0000_0888_3FE7
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a121_1 ( .OUT(na121_1_i), .IN1(~na3_1), .IN2(~na120_1), .IN3(na422_2), .IN4(na70_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(~na301_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a121_2 ( .OUT(na121_1), .CLK(~na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na121_1_i) );
// C_MX2a////      x12y42     80'h00_0018_00_0040_0C0A_4F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a122_1 ( .OUT(na122_1), .IN1(1'b0), .IN2(na8_1), .IN3(1'b0), .IN4(na113_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na53_2), .IN8(na107_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x11y40     80'h00_FE00_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a123_1 ( .OUT(na123_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na368_2), .IN6(na123_1), .IN7(na75_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a123_2 ( .OUT(na123_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na123_1_i) );
// C_ADDF2///ADDF2/      x9y39     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a126_1 ( .OUT(na126_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na4_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na148_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a126_4 ( .OUT(na126_2), .COUTY1(na126_4), .IN1(1'b0), .IN2(1'b0), .IN3(na4_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na148_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x9y40     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a128_1 ( .OUT(na128_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na100_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na126_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a128_4 ( .OUT(na128_2), .COUTY1(na128_4), .IN1(1'b1), .IN2(na100_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na100_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na126_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x9y41     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a130_1 ( .OUT(na130_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na36_2),
                     .CINX(1'b0), .CINY1(na128_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a130_4 ( .OUT(na130_2), .COUTY1(na130_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na36_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na36_2), .CINX(1'b0), .CINY1(na128_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x9y42     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a132_1 ( .OUT(na132_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na26_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na130_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a132_4 ( .OUT(na132_2), .COUTY1(na132_4), .IN1(1'b0), .IN2(1'b0), .IN3(na26_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na26_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na130_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x9y43     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a134_1 ( .OUT(na134_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na31_2),
                     .CINX(1'b0), .CINY1(na132_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a134_4 ( .OUT(na134_2), .COUTY1(na134_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na31_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na31_2), .CINX(1'b0), .CINY1(na132_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x9y34     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a135_1 ( .OUT(na135_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na62_2), .IN7(na42_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na149_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a135_4 ( .OUT(na135_2), .COUTY1(na135_4), .IN1(1'b1), .IN2(na62_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na62_2), .IN7(na42_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na149_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x9y44     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a137_1 ( .OUT(na137_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na27_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na134_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a137_4 ( .OUT(na137_2), .COUTY1(na137_4), .IN1(1'b1), .IN2(na27_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na27_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na134_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x9y45     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a139_1 ( .OUT(na139_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na13_2),
                     .CINX(1'b0), .CINY1(na137_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a139_4 ( .OUT(na139_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na13_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na13_2),
                     .CINX(1'b0), .CINY1(na137_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x9y35     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a142_1 ( .OUT(na142_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na40_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na135_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a142_4 ( .OUT(na142_2), .COUTY1(na142_4), .IN1(na40_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na40_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na135_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x9y36     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a144_1 ( .OUT(na144_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na63_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na142_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a144_4 ( .OUT(na144_2), .COUTY1(na144_4), .IN1(na63_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na63_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na142_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x9y37     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a146_1 ( .OUT(na146_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na37_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na144_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a146_4 ( .OUT(na146_2), .COUTY1(na146_4), .IN1(na37_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na37_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na144_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x9y38     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a148_1 ( .OUT(na148_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na47_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na146_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a148_4 ( .OUT(na148_2), .COUTY1(na148_4), .IN1(1'b1), .IN2(na47_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na47_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na146_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x9y33     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a149_2 ( .OUT(na149_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a149_6 ( .COUTY1(na149_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na149_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x19y38     80'h00_0078_00_0020_0C66_CCA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a150_1 ( .OUT(na150_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na88_1), .IN7(1'b1), .IN8(na87_1),
                     .CINX(1'b0), .CINY1(na158_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a150_4 ( .OUT(na150_2), .COUTY1(na150_4), .IN1(1'b0), .IN2(1'b0), .IN3(na89_1), .IN4(1'b1), .IN5(1'b1), .IN6(na88_1), .IN7(1'b1),
                     .IN8(na87_1), .CINX(1'b0), .CINY1(na158_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x19y39     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a152_1 ( .OUT(na152_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na90_1),
                     .CINX(1'b0), .CINY1(na150_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a152_4 ( .OUT(na152_2), .COUTY1(na152_4), .IN1(na91_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na90_1), .CINX(1'b0), .CINY1(na150_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x19y40     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a154_1 ( .OUT(na154_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na92_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na152_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a154_4 ( .OUT(na154_2), .COUTY1(na154_4), .IN1(na93_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na92_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na152_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x19y41     80'h00_0078_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a156_1 ( .OUT(na156_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na94_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na154_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a156_4 ( .OUT(na156_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na95_1), .IN5(1'b0), .IN6(1'b0), .IN7(na94_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na154_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x19y37     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a158_2 ( .OUT(na158_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a158_6 ( .COUTY1(na158_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na158_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x18y34     80'h00_0078_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a159_1 ( .OUT(na159_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na115_2), .IN7(na111_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na167_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a159_4 ( .OUT(na159_2), .COUTY1(na159_4), .IN1(1'b0), .IN2(1'b0), .IN3(na111_1), .IN4(1'b1), .IN5(1'b1), .IN6(na115_2), .IN7(na111_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na167_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x18y35     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a161_1 ( .OUT(na161_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na79_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na159_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a161_4 ( .OUT(na161_2), .COUTY1(na161_4), .IN1(na79_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na79_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na159_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x18y36     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a163_1 ( .OUT(na163_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na67_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na161_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a163_4 ( .OUT(na163_2), .COUTY1(na163_4), .IN1(1'b0), .IN2(1'b0), .IN3(na67_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na67_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na161_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x18y37     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a165_1 ( .OUT(na165_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na56_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na163_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a165_4 ( .OUT(na165_2), .IN1(na56_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na56_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na163_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x18y33     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a167_2 ( .OUT(na167_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a167_6 ( .COUTY1(na167_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na167_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x12y29     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a168_1 ( .OUT(na168_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na51_2), .IN6(1'b1), .IN7(1'b1), .IN8(na55_1),
                     .CINX(1'b0), .CINY1(na176_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a168_4 ( .OUT(na168_2), .COUTY1(na168_4), .IN1(na51_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na51_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na55_1), .CINX(1'b0), .CINY1(na176_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x12y30     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a170_1 ( .OUT(na170_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na49_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na168_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a170_4 ( .OUT(na170_2), .COUTY1(na170_4), .IN1(1'b1), .IN2(na49_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na49_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na168_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x12y31     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a172_1 ( .OUT(na172_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na17_2),
                     .CINX(1'b0), .CINY1(na170_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a172_4 ( .OUT(na172_2), .COUTY1(na172_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na38_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na17_2), .CINX(1'b0), .CINY1(na170_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x12y32     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a174_1 ( .OUT(na174_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na25_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na172_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a174_4 ( .OUT(na174_2), .IN1(1'b1), .IN2(na25_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na25_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na172_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x12y28     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a176_2 ( .OUT(na176_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a176_6 ( .COUTY1(na176_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na176_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x13y34     80'h00_0078_00_0020_0C66_ACC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a177_1 ( .OUT(na177_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na441_2), .IN7(na1_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na339_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a177_4 ( .OUT(na177_2), .COUTY1(na177_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na108_1), .IN5(1'b1), .IN6(na441_2), .IN7(na1_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na339_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x13y35     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a179_1 ( .OUT(na179_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na78_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na177_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a179_4 ( .OUT(na179_2), .COUTY1(na179_4), .IN1(1'b0), .IN2(1'b0), .IN3(na78_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na78_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na177_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x13y36     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a181_1 ( .OUT(na181_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na5_1),
                     .CINX(1'b0), .CINY1(na179_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a181_4 ( .OUT(na181_2), .COUTY1(na181_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na112_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na5_1), .CINX(1'b0), .CINY1(na179_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x13y37     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a183_1 ( .OUT(na183_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na106_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na181_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a183_4 ( .OUT(na183_2), .IN1(1'b0), .IN2(1'b0), .IN3(na43_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na106_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na181_4), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0014_0016)) 
           _a187 ( .GLB0(na187_1), .GLB1(na187_2), .GLB2(_d0), .GLB3(_d1), .CLK_FB0(_d2), .CLK_FB1(_d3), .CLK_FB2(_d4), .CLK_FB3(_d5),
                   .CLK0_0(na305_6), .CLK0_90(na305_5), .CLK0_180(na305_4), .CLK0_270(na305_3), .CLK0_BYP(1'b0), .CLK1_0(na304_6),
                   .CLK1_90(na304_5), .CLK1_180(na304_4), .CLK1_270(na304_3), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0),
                   .CLK2_270(1'b0), .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0),
                   .USR_GLB0(1'b0), .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0),
                   .USR_FB3(1'b0) );
// C_AND/D///      x17y43     80'h00_FE00_00_0000_0C88_F3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a204_1 ( .OUT(na204_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na20_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a204_2 ( .OUT(na204_1), .CLK(na300_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na204_1_i) );
// C_///AND/D      x12y44     80'h00_FE00_80_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a205_4 ( .OUT(na205_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na75_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a205_5 ( .OUT(na205_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na205_2_i) );
// C_AND/D///      x12y38     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a255_1 ( .OUT(na255_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na43_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a255_2 ( .OUT(na255_1), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na255_1_i) );
// C_///AND/D      x16y35     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a265_4 ( .OUT(na265_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na17_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a265_5 ( .OUT(na265_2), .CLK(na187_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na265_2_i) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a298 ( .Y(na298_1), .I(clk) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a299 ( .Y(na299_1), .I(i_mosi_ILA) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a300 ( .Y(na300_1), .I(i_sclk_ILA) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a301 ( .Y(na301_1), .I(i_ss_ILA) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a302 ( .O(led), .A(na369_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a303 ( .O(o_miso_ILA), .A(na370_10) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_0C_08_0C_20_82)) 
           _a304 ( .USR_PLL_LOCKED_STDY(_d6), .USR_PLL_LOCKED(_d7), .CLK270(na304_3), .CLK180(na304_4), .CLK90(na304_5), .CLK0(na304_6),
                   .CLK_REF_OUT(_d8), .CLK_REF(na308_2), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_73_08_17_10_82)) 
           _a305 ( .USR_PLL_LOCKED_STDY(_d9), .USR_PLL_LOCKED(_d10), .CLK270(na305_3), .CLK180(na305_4), .CLK90(na305_5), .CLK0(na305_6),
                   .CLK_REF_OUT(_d11), .CLK_REF(na308_1), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_01_04_05_00_60_00_0D_00_00_00_03_13_00_00_00_23_00_13_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a306 ( .DOA({_d12, _d13, _d14, _d15, _d16, _d17, _d18, _d19, _d20, _d21, _d22, _d23, _d24, _d25, _d26, _d27, _d28, _d29,
                  _d30, _d31, _d32, _d33, _d34, _d35, _d36, _d37, _d38, _d39, _d40, _d41, _d42, _d43, _d44, _d45, _d46, _d47, _d48,
                  _d49, _d50, _d51}),
                   .DOAX({_d52, _d53, _d54, _d55, _d56, _d57, _d58, _d59, _d60, _d61, _d62, _d63, _d64, _d65, _d66, _d67, _d68, _d69,
                  _d70, _d71, _d72, _d73, _d74, _d75, _d76, _d77, _d78, _d79, _d80, _d81, _d82, _d83, _d84, _d85, _d86, _d87, _d88,
                  _d89, _d90, _d91}),
                   .DOB({_d92, _d93, _d94, _d95, _d96, _d97, _d98, _d99, _d100, _d101, _d102, _d103, _d104, _d105, _d106, _d107, _d108,
                  _d109, _d110, _d111, _d112, _d113, _d114, _d115, _d116, _d117, _d118, _d119, _d120, _d121, _d122, _d123, _d124, _d125,
                  _d126, _d127, _d128, _d129, _d130, na306_120}),
                   .DOBX({_d131, _d132, _d133, _d134, _d135, _d136, _d137, _d138, _d139, _d140, _d141, _d142, _d143, _d144, _d145,
                  _d146, _d147, _d148, _d149, _d150, _d151, _d152, _d153, _d154, _d155, _d156, _d157, _d158, _d159, _d160, _d161, _d162,
                  _d163, _d164, _d165, _d166, _d167, _d168, _d169, _d170}),
                   .ECC1B_ERRA({_d171, _d172, _d173, _d174}),
                   .ECC1B_ERRB({_d175, _d176, _d177, _d178}),
                   .ECC2B_ERRA({_d179, _d180, _d181, _d182}),
                   .ECC2B_ERRB({_d183, _d184, _d185, _d186}),
                   .FORW_CAS_WRAO(_d187), .FORW_CAS_WRBO(_d188), .FORW_CAS_BMAO(_d189), .FORW_CAS_BMBO(_d190), .FORW_CAS_RDAO(_d191),
                   .FORW_CAS_RDBO(_d192), .FORW_UADDRAO({_d193, _d194, _d195, _d196, _d197, _d198, _d199, _d200, _d201, _d202, _d203,
                  _d204, _d205, _d206, _d207, _d208}),
                   .FORW_LADDRAO({_d209, _d210, _d211, _d212, _d213, _d214, _d215, _d216, _d217, _d218, _d219, _d220, _d221, _d222,
                  _d223, _d224}),
                   .FORW_UADDRBO({_d225, _d226, _d227, _d228, _d229, _d230, _d231, _d232, _d233, _d234, _d235, _d236, _d237, _d238,
                  _d239, _d240}),
                   .FORW_LADDRBO({_d241, _d242, _d243, _d244, _d245, _d246, _d247, _d248, _d249, _d250, _d251, _d252, _d253, _d254,
                  _d255, _d256}),
                   .FORW_UA0CLKO(_d257), .FORW_UA0ENO(_d258), .FORW_UA0WEO(_d259), .FORW_LA0CLKO(_d260), .FORW_LA0ENO(_d261), .FORW_LA0WEO(_d262),
                   .FORW_UA1CLKO(_d263), .FORW_UA1ENO(_d264), .FORW_UA1WEO(_d265), .FORW_LA1CLKO(_d266), .FORW_LA1ENO(_d267), .FORW_LA1WEO(_d268),
                   .FORW_UB0CLKO(_d269), .FORW_UB0ENO(_d270), .FORW_UB0WEO(_d271), .FORW_LB0CLKO(_d272), .FORW_LB0ENO(_d273), .FORW_LB0WEO(_d274),
                   .FORW_UB1CLKO(_d275), .FORW_UB1ENO(_d276), .FORW_UB1WEO(_d277), .FORW_LB1CLKO(_d278), .FORW_LB1ENO(_d279), .FORW_LB1WEO(_d280),
                   .CLOCKA({_d281, _d282, _d283, _d284}),
                   .CLOCKB({_d285, _d286, _d287, _d288}),
                   .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .CLKB({1'b1, 1'b1, 1'b1, na313_9}),
                   .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .GLWEA({1'b1, 1'b1, 1'b1, na314_10}),
                   .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0({na319_10, na326_9, na333_10, na336_9, na338_10, na340_9, na341_10, na342_9, na344_10, na345_9, na346_10,
                  na351_9, na353_10, na359_9, na360_10, na364_9}),
                   .ADDRA1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB0({na366_10, na367_9, na371_10, na372_9, na373_10, na374_9, na375_10, na376_9, na377_10, na378_9, na379_10,
                  na380_9, na381_10, na382_9, na383_10, na384_9}),
                   .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .DIA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, na385_10, na386_9, na387_10, na388_9, na389_10, na390_9, na391_10, na392_9, na393_10, na394_9, na395_10,
                  na396_9, na397_10, na398_9, na399_10, na400_9, na401_10, na402_9, na403_10, na404_9}),
                   .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, na405_10, na406_9, na407_10, na408_9, na409_10, na410_9, na411_10, na412_9, na413_10, na414_9, na415_10,
                  na416_9, na417_10, na418_9, na419_10, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .CLOCK1(na187_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                   .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                   .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                   .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                   .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
CC_USR_RSTN            _a307 ( .USR_RSTN(na307_1) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a308 ( .PCLK0(na308_1), .PCLK1(na308_2), .PCLK2(_d289), .PCLK3(_d290), .CLK0(na298_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0),
                   .SER_CLK(1'b0), .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_MX2b////      x12y37     80'h00_0018_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a309_1 ( .OUT(na309_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1_2), .IN4(1'b1), .IN5(1'b0), .IN6(na181_1), .IN7(1'b0), .IN8(na5_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x16y35     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a310_1 ( .OUT(na310_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na24_1), .IN6(1'b1), .IN7(1'b1), .IN8(na428_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x11y38     80'h00_0018_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a311_1 ( .OUT(na311_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1_2), .IN4(1'b1), .IN5(na179_1), .IN6(1'b0), .IN7(na78_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x1y66     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a312_5 ( .OUT(na312_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na307_1), .CP_O(1'b0) );
// C_AND////      x35y33     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a313_1 ( .OUT(na313_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na300_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a313_6 ( .RAM_O1(na313_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na313_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x27y33     80'h08_0060_00_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a314_4 ( .OUT(na314_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na55_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a314_6 ( .RAM_O2(na314_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na314_2), .COMP_OUT(1'b0) );
// C_MX2b////      x22y31     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a315_1 ( .OUT(na315_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na55_2), .IN5(1'b0), .IN6(na25_1), .IN7(1'b0), .IN8(na174_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x14y30     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a316_1 ( .OUT(na316_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na55_2), .IN5(1'b0), .IN6(na25_2), .IN7(1'b0), .IN8(na174_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x20y38     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a317_1 ( .OUT(na317_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na32_1), .IN7(1'b0), .IN8(na429_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x17y31     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a318_1 ( .OUT(na318_1), .IN1(1'b1), .IN2(na433_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na172_2), .IN8(na38_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a319_4 ( .OUT(na319_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a319_6 ( .RAM_O2(na319_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na319_2), .COMP_OUT(1'b0) );
// C_MX2b////      x16y27     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a320_1 ( .OUT(na320_1), .IN1(1'b1), .IN2(na433_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na172_1), .IN8(na17_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x14y29     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a321_1 ( .OUT(na321_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na55_2), .IN5(1'b0), .IN6(na49_1), .IN7(1'b0), .IN8(na170_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x18y29     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a322_1 ( .OUT(na322_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na55_2), .IN5(1'b0), .IN6(na49_2), .IN7(1'b0), .IN8(na170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x16y29     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a323_1 ( .OUT(na323_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na55_2), .IN5(na51_1), .IN6(1'b0), .IN7(na168_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x15y28     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a324_1 ( .OUT(na324_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na55_2), .IN5(na51_2), .IN6(1'b0), .IN7(na168_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x14y42     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a325_1 ( .OUT(na325_1), .IN1(1'b1), .IN2(na54_2), .IN3(1'b0), .IN4(1'b0), .IN5(na431_2), .IN6(na2_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a326_1 ( .OUT(na326_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a326_6 ( .RAM_O1(na326_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na326_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x17y30     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a327_1 ( .OUT(na327_1), .IN1(1'b1), .IN2(~na433_2), .IN3(1'b0), .IN4(1'b0), .IN5(na56_1), .IN6(na25_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x16y31     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a328_1 ( .OUT(na328_1), .IN1(1'b1), .IN2(~na433_2), .IN3(1'b0), .IN4(1'b0), .IN5(na56_2), .IN6(na25_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x17y41     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a329_1 ( .OUT(na329_1), .IN1(na59_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na58_1), .IN8(na33_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x16y43     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a330_1 ( .OUT(na330_1), .IN1(na59_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na434_2), .IN6(na2_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x24y31     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a331_1 ( .OUT(na331_1), .IN1(1'b1), .IN2(~na433_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na67_1), .IN8(na38_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x21y34     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a332_1 ( .OUT(na332_1), .IN1(1'b1), .IN2(~na433_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na67_2), .IN8(na17_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a333_4 ( .OUT(na333_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a333_6 ( .RAM_O2(na333_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na333_2), .COMP_OUT(1'b0) );
// C_///AND/      x24y37     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a334_4 ( .OUT(na334_2), .IN1(1'b1), .IN2(na110_1), .IN3(1'b1), .IN4(na429_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x22y36     80'h00_0018_00_0000_0888_C5DC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a335_1 ( .OUT(na335_1), .IN1(1'b0), .IN2(na437_2), .IN3(~na424_2), .IN4(na55_2), .IN5(~na446_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na73_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y39     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a336_1 ( .OUT(na336_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na56_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a336_6 ( .RAM_O1(na336_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na336_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x16y33     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a337_4 ( .OUT(na337_2), .IN1(~na24_2), .IN2(1'b1), .IN3(1'b1), .IN4(na55_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y38     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a338_4 ( .OUT(na338_2), .IN1(na56_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a338_6 ( .RAM_O2(na338_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na338_2), .COMP_OUT(1'b0) );
// C_/C_0_1///      x13y33     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a339_2 ( .OUT(na339_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a339_6 ( .COUTY1(na339_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na339_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x28y38     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a340_1 ( .OUT(na340_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na67_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a340_6 ( .RAM_O1(na340_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na340_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y37     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a341_4 ( .OUT(na341_2), .IN1(1'b1), .IN2(1'b1), .IN3(na67_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a341_6 ( .RAM_O2(na341_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na341_2), .COMP_OUT(1'b0) );
// C_AND////      x28y37     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a342_1 ( .OUT(na342_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na79_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a342_6 ( .RAM_O1(na342_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na342_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x18y32     80'h00_0018_00_0000_0888_C5DC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a343_1 ( .OUT(na343_1), .IN1(1'b0), .IN2(na437_2), .IN3(~na16_2), .IN4(na55_2), .IN5(~na446_2), .IN6(1'b0), .IN7(1'b0), .IN8(na73_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y36     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a344_4 ( .OUT(na344_2), .IN1(na79_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a344_6 ( .RAM_O2(na344_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na344_2), .COMP_OUT(1'b0) );
// C_AND////      x28y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a345_1 ( .OUT(na345_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a345_6 ( .RAM_O1(na345_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na345_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y35     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a346_4 ( .OUT(na346_2), .IN1(1'b1), .IN2(1'b1), .IN3(na111_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a346_6 ( .RAM_O2(na346_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na346_2), .COMP_OUT(1'b0) );
// C_MX2b////      x12y34     80'h00_0018_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a347_1 ( .OUT(na347_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1_2), .IN4(1'b1), .IN5(na179_2), .IN6(1'b0), .IN7(na78_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x19y33     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a348_1 ( .OUT(na348_1), .IN1(1'b1), .IN2(~na433_2), .IN3(1'b0), .IN4(1'b0), .IN5(na79_1), .IN6(na49_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x24y35     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a349_1 ( .OUT(na349_1), .IN1(1'b1), .IN2(~na433_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na111_2), .IN8(na55_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x14y38     80'h00_0018_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a350_1 ( .OUT(na350_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1_2), .IN4(1'b1), .IN5(1'b0), .IN6(na177_1), .IN7(1'b0), .IN8(na108_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y35     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a351_1 ( .OUT(na351_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na115_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a351_6 ( .RAM_O1(na351_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na351_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x16y30     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a352_1 ( .OUT(na352_1), .IN1(1'b1), .IN2(~na433_2), .IN3(1'b0), .IN4(1'b0), .IN5(na79_2), .IN6(na49_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y34     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a353_4 ( .OUT(na353_2), .IN1(1'b1), .IN2(1'b1), .IN3(na111_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a353_6 ( .RAM_O2(na353_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na353_2), .COMP_OUT(1'b0) );
// C_MX2b////      x16y46     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a354_1 ( .OUT(na354_1), .IN1(~na59_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na61_1), .IN8(na440_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x10y38     80'h00_0018_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a355_1 ( .OUT(na355_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1_2), .IN4(1'b1), .IN5(na183_2), .IN6(1'b0), .IN7(na43_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x15y38     80'h00_0018_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a356_1 ( .OUT(na356_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1_2), .IN4(1'b1), .IN5(na183_1), .IN6(1'b0), .IN7(na106_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x14y43     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a357_1 ( .OUT(na357_1), .IN1(1'b1), .IN2(~na54_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na61_1), .IN8(na107_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x13y32     80'h00_0018_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a358_1 ( .OUT(na358_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1_2), .IN4(1'b1), .IN5(1'b0), .IN6(na177_2), .IN7(1'b0), .IN8(na108_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a359_1 ( .OUT(na359_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a359_6 ( .RAM_O1(na359_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na359_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a360_4 ( .OUT(na360_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a360_6 ( .RAM_O2(na360_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na360_2), .COMP_OUT(1'b0) );
// C_MX2b////      x22y37     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a361_1 ( .OUT(na361_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na55_2), .IN5(na51_1), .IN6(1'b0), .IN7(na111_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x14y40     80'h00_0018_00_0040_0AA0_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a362_1 ( .OUT(na362_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1_2), .IN4(1'b1), .IN5(1'b0), .IN6(na181_2), .IN7(1'b0), .IN8(na112_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x20y30     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a363_1 ( .OUT(na363_1), .IN1(1'b1), .IN2(na433_2), .IN3(1'b0), .IN4(1'b0), .IN5(na51_2), .IN6(na115_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a364_1 ( .OUT(na364_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a364_6 ( .RAM_O1(na364_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na364_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x24y38     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a365_1 ( .OUT(na365_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na24_2), .IN6(na110_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a366_4 ( .OUT(na366_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a366_6 ( .RAM_O2(na366_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na366_2), .COMP_OUT(1'b0) );
// C_AND////      x37y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a367_1 ( .OUT(na367_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a367_6 ( .RAM_O1(na367_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na367_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x13y39     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a368_4 ( .OUT(na368_2), .IN1(na109_1), .IN2(1'b1), .IN3(1'b1), .IN4(na122_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x1y95     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a369_4 ( .OUT(na369_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na13_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a369_6 ( .RAM_O2(na369_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na369_2), .COMP_OUT(1'b0) );
// C_///AND/      x19y1     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a370_4 ( .OUT(na370_2), .IN1(na76_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a370_6 ( .RAM_O2(na370_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na370_2), .COMP_OUT(1'b0) );
// C_///AND/      x37y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a371_4 ( .OUT(na371_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a371_6 ( .RAM_O2(na371_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na371_2), .COMP_OUT(1'b0) );
// C_AND////      x37y39     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a372_1 ( .OUT(na372_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na95_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a372_6 ( .RAM_O1(na372_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na372_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y38     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a373_4 ( .OUT(na373_2), .IN1(1'b1), .IN2(1'b1), .IN3(na94_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a373_6 ( .RAM_O2(na373_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na373_2), .COMP_OUT(1'b0) );
// C_AND////      x37y38     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a374_1 ( .OUT(na374_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na93_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a374_6 ( .RAM_O1(na374_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na374_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y37     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a375_4 ( .OUT(na375_2), .IN1(1'b1), .IN2(1'b1), .IN3(na92_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a375_6 ( .RAM_O2(na375_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na375_2), .COMP_OUT(1'b0) );
// C_AND////      x37y37     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a376_1 ( .OUT(na376_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na91_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a376_6 ( .RAM_O1(na376_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na376_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y36     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a377_4 ( .OUT(na377_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na90_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a377_6 ( .RAM_O2(na377_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na377_2), .COMP_OUT(1'b0) );
// C_AND////      x37y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a378_1 ( .OUT(na378_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a378_6 ( .RAM_O1(na378_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na378_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y35     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a379_4 ( .OUT(na379_2), .IN1(1'b1), .IN2(1'b1), .IN3(na89_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a379_6 ( .RAM_O2(na379_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na379_2), .COMP_OUT(1'b0) );
// C_AND////      x37y35     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a380_1 ( .OUT(na380_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na88_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a380_6 ( .RAM_O1(na380_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na380_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y34     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a381_4 ( .OUT(na381_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na87_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a381_6 ( .RAM_O2(na381_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na381_2), .COMP_OUT(1'b0) );
// C_AND////      x37y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a382_1 ( .OUT(na382_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a382_6 ( .RAM_O1(na382_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na382_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a383_4 ( .OUT(na383_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a383_6 ( .RAM_O2(na383_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na383_2), .COMP_OUT(1'b0) );
// C_AND////      x37y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a384_1 ( .OUT(na384_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a384_6 ( .RAM_O1(na384_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na384_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a385_4 ( .OUT(na385_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a385_6 ( .RAM_O2(na385_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na385_2), .COMP_OUT(1'b0) );
// C_AND////      x30y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a386_1 ( .OUT(na386_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a386_6 ( .RAM_O1(na386_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na386_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a387_4 ( .OUT(na387_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a387_6 ( .RAM_O2(na387_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na387_2), .COMP_OUT(1'b0) );
// C_AND////      x30y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a388_1 ( .OUT(na388_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a388_6 ( .RAM_O1(na388_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na388_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a389_4 ( .OUT(na389_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a389_6 ( .RAM_O2(na389_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na389_2), .COMP_OUT(1'b0) );
// C_AND////      x32y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a390_1 ( .OUT(na390_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a390_6 ( .RAM_O1(na390_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na390_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a391_4 ( .OUT(na391_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a391_6 ( .RAM_O2(na391_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na391_2), .COMP_OUT(1'b0) );
// C_AND////      x32y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a392_1 ( .OUT(na392_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a392_6 ( .RAM_O1(na392_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na392_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y38     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a393_4 ( .OUT(na393_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a393_6 ( .RAM_O2(na393_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na393_2), .COMP_OUT(1'b0) );
// C_AND////      x32y38     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a394_1 ( .OUT(na394_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a394_6 ( .RAM_O1(na394_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na394_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y37     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a395_4 ( .OUT(na395_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a395_6 ( .RAM_O2(na395_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na395_2), .COMP_OUT(1'b0) );
// C_AND////      x32y37     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a396_1 ( .OUT(na396_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a396_6 ( .RAM_O1(na396_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na396_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y36     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a397_4 ( .OUT(na397_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a397_6 ( .RAM_O2(na397_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na397_2), .COMP_OUT(1'b0) );
// C_AND////      x32y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a398_1 ( .OUT(na398_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a398_6 ( .RAM_O1(na398_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na398_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y35     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a399_4 ( .OUT(na399_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a399_6 ( .RAM_O2(na399_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na399_2), .COMP_OUT(1'b0) );
// C_AND////      x32y35     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a400_1 ( .OUT(na400_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a400_6 ( .RAM_O1(na400_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na400_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y34     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a401_4 ( .OUT(na401_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a401_6 ( .RAM_O2(na401_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na401_2), .COMP_OUT(1'b0) );
// C_AND////      x32y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a402_1 ( .OUT(na402_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a402_6 ( .RAM_O1(na402_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na402_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a403_4 ( .OUT(na403_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a403_6 ( .RAM_O2(na403_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na403_2), .COMP_OUT(1'b0) );
// C_AND////      x32y33     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a404_1 ( .OUT(na404_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na298_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a404_6 ( .RAM_O1(na404_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na404_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a405_4 ( .OUT(na405_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a405_6 ( .RAM_O2(na405_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na405_2), .COMP_OUT(1'b0) );
// C_AND////      x29y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a406_1 ( .OUT(na406_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a406_6 ( .RAM_O1(na406_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na406_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a407_4 ( .OUT(na407_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a407_6 ( .RAM_O2(na407_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na407_2), .COMP_OUT(1'b0) );
// C_AND////      x29y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a408_1 ( .OUT(na408_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a408_6 ( .RAM_O1(na408_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na408_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a409_4 ( .OUT(na409_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a409_6 ( .RAM_O2(na409_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na409_2), .COMP_OUT(1'b0) );
// C_AND////      x31y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a410_1 ( .OUT(na410_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a410_6 ( .RAM_O1(na410_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na410_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a411_4 ( .OUT(na411_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a411_6 ( .RAM_O2(na411_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na411_2), .COMP_OUT(1'b0) );
// C_AND////      x31y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a412_1 ( .OUT(na412_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a412_6 ( .RAM_O1(na412_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na412_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y38     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a413_4 ( .OUT(na413_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a413_6 ( .RAM_O2(na413_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na413_2), .COMP_OUT(1'b0) );
// C_AND////      x31y38     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a414_1 ( .OUT(na414_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a414_6 ( .RAM_O1(na414_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na414_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y37     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a415_4 ( .OUT(na415_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a415_6 ( .RAM_O2(na415_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na415_2), .COMP_OUT(1'b0) );
// C_AND////      x31y37     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a416_1 ( .OUT(na416_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a416_6 ( .RAM_O1(na416_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na416_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y36     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a417_4 ( .OUT(na417_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a417_6 ( .RAM_O2(na417_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na417_2), .COMP_OUT(1'b0) );
// C_AND////      x31y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a418_1 ( .OUT(na418_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a418_6 ( .RAM_O1(na418_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na418_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y35     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a419_4 ( .OUT(na419_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a419_6 ( .RAM_O2(na419_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na419_2), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x34y33     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a420_2 ( .OUT(na420_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na306_120), .CP_O(1'b0) );
// C_////Bridge      x14y36     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a421_5 ( .OUT(na421_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1_1), .IN8(1'b0) );
// C_////Bridge      x22y31     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a422_5 ( .OUT(na422_2), .IN1(na3_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x18y42     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a423_5 ( .OUT(na423_2), .IN1(na9_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y35     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a424_5 ( .OUT(na424_2), .IN1(na9_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y42     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a425_5 ( .OUT(na425_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na16_2), .IN8(1'b0) );
// C_////Bridge      x18y33     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a426_5 ( .OUT(na426_2), .IN1(1'b0), .IN2(na20_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x14y30     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a427_5 ( .OUT(na427_2), .IN1(1'b0), .IN2(na20_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y38     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a428_5 ( .OUT(na428_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na24_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x16y36     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a429_5 ( .OUT(na429_2), .IN1(1'b0), .IN2(na34_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x16y40     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a430_5 ( .OUT(na430_2), .IN1(na44_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x11y39     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a431_5 ( .OUT(na431_2), .IN1(1'b0), .IN2(1'b0), .IN3(na53_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x18y31     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a432_5 ( .OUT(na432_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na55_1) );
// C_////Bridge      x19y30     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a433_5 ( .OUT(na433_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na55_2) );
// C_////Bridge      x17y43     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a434_5 ( .OUT(na434_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na60_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y34     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a435_5 ( .OUT(na435_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na73_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y37     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a436_5 ( .OUT(na436_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na73_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y34     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a437_5 ( .OUT(na437_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na73_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y46     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a438_5 ( .OUT(na438_2), .IN1(1'b0), .IN2(1'b0), .IN3(na75_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y45     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a439_5 ( .OUT(na439_2), .IN1(1'b0), .IN2(na101_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x18y46     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a440_5 ( .OUT(na440_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na104_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x13y32     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a441_5 ( .OUT(na441_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na108_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x18y32     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a442_5 ( .OUT(na442_2), .IN1(na109_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x12y34     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a443_5 ( .OUT(na443_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na123_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x10y45     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a444_5 ( .OUT(na444_2), .IN1(1'b0), .IN2(na312_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x11y43     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a445_5 ( .OUT(na445_2), .IN1(1'b0), .IN2(na312_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y33     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a446_5 ( .OUT(na446_2), .IN1(1'b0), .IN2(1'b0), .IN3(na337_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
endmodule
