
module progmem (
    // Clock & reset
    input wire clk,
    input wire rstn,

    // PicoRV32 bus interface
    input  wire        valid,
    output wire        ready,	
    input  wire [31:0] addr,
    output wire [31:0] rdata,
	// Rewrite firmware
    input  wire        wen,
	input  wire [31:0] waddr,
	input  wire [31:0] wdata
);

  // ============================================================================

  localparam MEM_SIZE_BITS = 13;  // In 32-bit words
  localparam MEM_SIZE = 1 << MEM_SIZE_BITS;
  localparam MEM_ADDR_MASK = 32'h0010_0000;

  // ============================================================================

  wire [MEM_SIZE_BITS-1:0] mem_addr;
  reg  [             31:0] mem_data;
  reg  [             31:0] mem      [0:MEM_SIZE];

  initial begin
    mem['h0000] <= 32'h00000093;
    mem['h0001] <= 32'h00000193;
    mem['h0002] <= 32'h00000213;
    mem['h0003] <= 32'h00000293;
    mem['h0004] <= 32'h00000313;
    mem['h0005] <= 32'h00000393;
    mem['h0006] <= 32'h00000413;
    mem['h0007] <= 32'h00000493;
    mem['h0008] <= 32'h00000513;
    mem['h0009] <= 32'h00000593;
    mem['h000A] <= 32'h00000613;
    mem['h000B] <= 32'h00000693;
    mem['h000C] <= 32'h00000713;
    mem['h000D] <= 32'h00000793;
    mem['h000E] <= 32'h00000813;
    mem['h000F] <= 32'h00000893;
    mem['h0010] <= 32'h00000913;
    mem['h0011] <= 32'h00000993;
    mem['h0012] <= 32'h00000A13;
    mem['h0013] <= 32'h00000A93;
    mem['h0014] <= 32'h00000B13;
    mem['h0015] <= 32'h00000B93;
    mem['h0016] <= 32'h00000C13;
    mem['h0017] <= 32'h00000C93;
    mem['h0018] <= 32'h00000D13;
    mem['h0019] <= 32'h00000D93;
    mem['h001A] <= 32'h00000E13;
    mem['h001B] <= 32'h00000E93;
    mem['h001C] <= 32'h00000F13;
    mem['h001D] <= 32'h00000F93;
    mem['h001E] <= 32'h00000513;
    mem['h001F] <= 32'h00000593;
    mem['h0020] <= 32'h00B52023;
    mem['h0021] <= 32'h00450513;
    mem['h0022] <= 32'hFE254CE3;
    mem['h0023] <= 32'h00005517;
    mem['h0024] <= 32'h47850513;
    mem['h0025] <= 32'h00000593;
    mem['h0026] <= 32'h07C00613;
    mem['h0027] <= 32'h00C5DC63;
    mem['h0028] <= 32'h00052683;
    mem['h0029] <= 32'h00D5A023;
    mem['h002A] <= 32'h00450513;
    mem['h002B] <= 32'h00458593;
    mem['h002C] <= 32'hFEC5C8E3;
    mem['h002D] <= 32'h07C00513;
    mem['h002E] <= 32'h53000593;
    mem['h002F] <= 32'h00B55863;
    mem['h0030] <= 32'h00052023;
    mem['h0031] <= 32'h00450513;
    mem['h0032] <= 32'hFEB54CE3;
    mem['h0033] <= 32'h534040EF;
    mem['h0034] <= 32'h0000006F;
    mem['h0035] <= 32'hFF010113;
    mem['h0036] <= 32'h00812623;
    mem['h0037] <= 32'h01010413;
    mem['h0038] <= 32'h030007B7;
    mem['h0039] <= 32'h0007A783;
    mem['h003A] <= 32'h0107D793;
    mem['h003B] <= 32'h0FF7F713;
    mem['h003C] <= 32'h52E00623;
    mem['h003D] <= 32'h00000013;
    mem['h003E] <= 32'h00C12403;
    mem['h003F] <= 32'h01010113;
    mem['h0040] <= 32'h00008067;
    mem['h0041] <= 32'hFE010113;
    mem['h0042] <= 32'h00812E23;
    mem['h0043] <= 32'h02010413;
    mem['h0044] <= 32'h00300793;
    mem['h0045] <= 32'hFEF406A3;
    mem['h0046] <= 32'hFE0407A3;
    mem['h0047] <= 32'h4A80006F;
    mem['h0048] <= 32'hFE040723;
    mem['h0049] <= 32'h4880006F;
    mem['h004A] <= 32'hFEF44703;
    mem['h004B] <= 32'h00070793;
    mem['h004C] <= 32'h00279793;
    mem['h004D] <= 32'h00E787B3;
    mem['h004E] <= 32'h00379793;
    mem['h004F] <= 32'h00078713;
    mem['h0050] <= 32'hFEE44783;
    mem['h0051] <= 32'h00F707B3;
    mem['h0052] <= 32'h00279713;
    mem['h0053] <= 32'h052007B7;
    mem['h0054] <= 32'h00F707B3;
    mem['h0055] <= 32'h00900713;
    mem['h0056] <= 32'h00E7A023;
    mem['h0057] <= 32'hFEF44703;
    mem['h0058] <= 32'hFED44783;
    mem['h0059] <= 32'h00F70A63;
    mem['h005A] <= 32'hFEF44703;
    mem['h005B] <= 32'hFED44783;
    mem['h005C] <= 32'h00478793;
    mem['h005D] <= 32'h00F71E63;
    mem['h005E] <= 32'hFEE44703;
    mem['h005F] <= 32'h00500793;
    mem['h0060] <= 32'h00E7F863;
    mem['h0061] <= 32'hFEE44703;
    mem['h0062] <= 32'h00800793;
    mem['h0063] <= 32'h02E7FC63;
    mem['h0064] <= 32'hFEE44703;
    mem['h0065] <= 32'h00600793;
    mem['h0066] <= 32'h00F70863;
    mem['h0067] <= 32'hFEE44703;
    mem['h0068] <= 32'h00800793;
    mem['h0069] <= 32'h04F71A63;
    mem['h006A] <= 32'hFEF44703;
    mem['h006B] <= 32'hFED44783;
    mem['h006C] <= 32'h04F76463;
    mem['h006D] <= 32'hFEF44703;
    mem['h006E] <= 32'hFED44783;
    mem['h006F] <= 32'h00478793;
    mem['h0070] <= 32'h02E7CC63;
    mem['h0071] <= 32'hFEF44703;
    mem['h0072] <= 32'h00070793;
    mem['h0073] <= 32'h00279793;
    mem['h0074] <= 32'h00E787B3;
    mem['h0075] <= 32'h00379793;
    mem['h0076] <= 32'h00078713;
    mem['h0077] <= 32'hFEE44783;
    mem['h0078] <= 32'h00F707B3;
    mem['h0079] <= 32'h00279713;
    mem['h007A] <= 32'h052007B7;
    mem['h007B] <= 32'h00F707B3;
    mem['h007C] <= 32'h00100713;
    mem['h007D] <= 32'h00E7A023;
    mem['h007E] <= 32'hFEF44703;
    mem['h007F] <= 32'hFED44783;
    mem['h0080] <= 32'h00F70A63;
    mem['h0081] <= 32'hFEF44703;
    mem['h0082] <= 32'hFED44783;
    mem['h0083] <= 32'h00278793;
    mem['h0084] <= 32'h00F71E63;
    mem['h0085] <= 32'hFEE44703;
    mem['h0086] <= 32'h00900793;
    mem['h0087] <= 32'h00E7F863;
    mem['h0088] <= 32'hFEE44703;
    mem['h0089] <= 32'h00C00793;
    mem['h008A] <= 32'h04E7FA63;
    mem['h008B] <= 32'hFEE44703;
    mem['h008C] <= 32'h00A00793;
    mem['h008D] <= 32'h02F71063;
    mem['h008E] <= 32'hFEF44703;
    mem['h008F] <= 32'hFED44783;
    mem['h0090] <= 32'h00F76A63;
    mem['h0091] <= 32'hFEF44703;
    mem['h0092] <= 32'hFED44783;
    mem['h0093] <= 32'h00478793;
    mem['h0094] <= 32'h02E7D663;
    mem['h0095] <= 32'hFEE44703;
    mem['h0096] <= 32'h00C00793;
    mem['h0097] <= 32'h04F71A63;
    mem['h0098] <= 32'hFEF44703;
    mem['h0099] <= 32'hFED44783;
    mem['h009A] <= 32'h04F76463;
    mem['h009B] <= 32'hFEF44703;
    mem['h009C] <= 32'hFED44783;
    mem['h009D] <= 32'h00278793;
    mem['h009E] <= 32'h02E7CC63;
    mem['h009F] <= 32'hFEF44703;
    mem['h00A0] <= 32'h00070793;
    mem['h00A1] <= 32'h00279793;
    mem['h00A2] <= 32'h00E787B3;
    mem['h00A3] <= 32'h00379793;
    mem['h00A4] <= 32'h00078713;
    mem['h00A5] <= 32'hFEE44783;
    mem['h00A6] <= 32'h00F707B3;
    mem['h00A7] <= 32'h00279713;
    mem['h00A8] <= 32'h052007B7;
    mem['h00A9] <= 32'h00F707B3;
    mem['h00AA] <= 32'h00100713;
    mem['h00AB] <= 32'h00E7A023;
    mem['h00AC] <= 32'hFEF44703;
    mem['h00AD] <= 32'hFED44783;
    mem['h00AE] <= 32'h02F70263;
    mem['h00AF] <= 32'hFEF44703;
    mem['h00B0] <= 32'hFED44783;
    mem['h00B1] <= 32'h00278793;
    mem['h00B2] <= 32'h00F70A63;
    mem['h00B3] <= 32'hFEF44703;
    mem['h00B4] <= 32'hFED44783;
    mem['h00B5] <= 32'h00478793;
    mem['h00B6] <= 32'h00F71E63;
    mem['h00B7] <= 32'hFEE44703;
    mem['h00B8] <= 32'h00D00793;
    mem['h00B9] <= 32'h00E7F863;
    mem['h00BA] <= 32'hFEE44703;
    mem['h00BB] <= 32'h01000793;
    mem['h00BC] <= 32'h02E7F663;
    mem['h00BD] <= 32'hFEE44703;
    mem['h00BE] <= 32'h00E00793;
    mem['h00BF] <= 32'h04F71A63;
    mem['h00C0] <= 32'hFEF44703;
    mem['h00C1] <= 32'hFED44783;
    mem['h00C2] <= 32'h04F76463;
    mem['h00C3] <= 32'hFEF44703;
    mem['h00C4] <= 32'hFED44783;
    mem['h00C5] <= 32'h00478793;
    mem['h00C6] <= 32'h02E7CC63;
    mem['h00C7] <= 32'hFEF44703;
    mem['h00C8] <= 32'h00070793;
    mem['h00C9] <= 32'h00279793;
    mem['h00CA] <= 32'h00E787B3;
    mem['h00CB] <= 32'h00379793;
    mem['h00CC] <= 32'h00078713;
    mem['h00CD] <= 32'hFEE44783;
    mem['h00CE] <= 32'h00F707B3;
    mem['h00CF] <= 32'h00279713;
    mem['h00D0] <= 32'h052007B7;
    mem['h00D1] <= 32'h00F707B3;
    mem['h00D2] <= 32'h00100713;
    mem['h00D3] <= 32'h00E7A023;
    mem['h00D4] <= 32'hFEF44703;
    mem['h00D5] <= 32'hFED44783;
    mem['h00D6] <= 32'h00F71E63;
    mem['h00D7] <= 32'hFEE44703;
    mem['h00D8] <= 32'h01100793;
    mem['h00D9] <= 32'h00E7F863;
    mem['h00DA] <= 32'hFEE44703;
    mem['h00DB] <= 32'h01400793;
    mem['h00DC] <= 32'h02E7FC63;
    mem['h00DD] <= 32'hFEE44703;
    mem['h00DE] <= 32'h01200793;
    mem['h00DF] <= 32'h00F70863;
    mem['h00E0] <= 32'hFEE44703;
    mem['h00E1] <= 32'h01400793;
    mem['h00E2] <= 32'h04F71A63;
    mem['h00E3] <= 32'hFEF44703;
    mem['h00E4] <= 32'hFED44783;
    mem['h00E5] <= 32'h04F76463;
    mem['h00E6] <= 32'hFEF44703;
    mem['h00E7] <= 32'hFED44783;
    mem['h00E8] <= 32'h00478793;
    mem['h00E9] <= 32'h02E7CC63;
    mem['h00EA] <= 32'hFEF44703;
    mem['h00EB] <= 32'h00070793;
    mem['h00EC] <= 32'h00279793;
    mem['h00ED] <= 32'h00E787B3;
    mem['h00EE] <= 32'h00379793;
    mem['h00EF] <= 32'h00078713;
    mem['h00F0] <= 32'hFEE44783;
    mem['h00F1] <= 32'h00F707B3;
    mem['h00F2] <= 32'h00279713;
    mem['h00F3] <= 32'h052007B7;
    mem['h00F4] <= 32'h00F707B3;
    mem['h00F5] <= 32'h00100713;
    mem['h00F6] <= 32'h00E7A023;
    mem['h00F7] <= 32'hFEE44703;
    mem['h00F8] <= 32'h01600793;
    mem['h00F9] <= 32'h00F70863;
    mem['h00FA] <= 32'hFEE44703;
    mem['h00FB] <= 32'h01800793;
    mem['h00FC] <= 32'h02F71863;
    mem['h00FD] <= 32'hFEF44703;
    mem['h00FE] <= 32'hFED44783;
    mem['h00FF] <= 32'h02F76263;
    mem['h0100] <= 32'hFEF44703;
    mem['h0101] <= 32'hFED44783;
    mem['h0102] <= 32'h00478793;
    mem['h0103] <= 32'h00E7CA63;
    mem['h0104] <= 32'hFEF44703;
    mem['h0105] <= 32'hFED44783;
    mem['h0106] <= 32'h00278793;
    mem['h0107] <= 32'h02F71063;
    mem['h0108] <= 32'hFEE44703;
    mem['h0109] <= 32'h01700793;
    mem['h010A] <= 32'h04F71463;
    mem['h010B] <= 32'hFEF44703;
    mem['h010C] <= 32'hFED44783;
    mem['h010D] <= 32'h00278793;
    mem['h010E] <= 32'h02F71C63;
    mem['h010F] <= 32'hFEF44703;
    mem['h0110] <= 32'h00070793;
    mem['h0111] <= 32'h00279793;
    mem['h0112] <= 32'h00E787B3;
    mem['h0113] <= 32'h00379793;
    mem['h0114] <= 32'h00078713;
    mem['h0115] <= 32'hFEE44783;
    mem['h0116] <= 32'h00F707B3;
    mem['h0117] <= 32'h00279713;
    mem['h0118] <= 32'h052007B7;
    mem['h0119] <= 32'h00F707B3;
    mem['h011A] <= 32'h00200713;
    mem['h011B] <= 32'h00E7A023;
    mem['h011C] <= 32'hFEF44703;
    mem['h011D] <= 32'hFED44783;
    mem['h011E] <= 32'h00F70A63;
    mem['h011F] <= 32'hFEF44703;
    mem['h0120] <= 32'hFED44783;
    mem['h0121] <= 32'h00478793;
    mem['h0122] <= 32'h00F71E63;
    mem['h0123] <= 32'hFEE44703;
    mem['h0124] <= 32'h01900793;
    mem['h0125] <= 32'h00E7F863;
    mem['h0126] <= 32'hFEE44703;
    mem['h0127] <= 32'h01C00793;
    mem['h0128] <= 32'h02E7F663;
    mem['h0129] <= 32'hFEE44703;
    mem['h012A] <= 32'h01A00793;
    mem['h012B] <= 32'h04F71A63;
    mem['h012C] <= 32'hFEF44703;
    mem['h012D] <= 32'hFED44783;
    mem['h012E] <= 32'h04F76463;
    mem['h012F] <= 32'hFEF44703;
    mem['h0130] <= 32'hFED44783;
    mem['h0131] <= 32'h00478793;
    mem['h0132] <= 32'h02E7CC63;
    mem['h0133] <= 32'hFEF44703;
    mem['h0134] <= 32'h00070793;
    mem['h0135] <= 32'h00279793;
    mem['h0136] <= 32'h00E787B3;
    mem['h0137] <= 32'h00379793;
    mem['h0138] <= 32'h00078713;
    mem['h0139] <= 32'hFEE44783;
    mem['h013A] <= 32'h00F707B3;
    mem['h013B] <= 32'h00279713;
    mem['h013C] <= 32'h052007B7;
    mem['h013D] <= 32'h00F707B3;
    mem['h013E] <= 32'h00200713;
    mem['h013F] <= 32'h00E7A023;
    mem['h0140] <= 32'hFEF44703;
    mem['h0141] <= 32'hFED44783;
    mem['h0142] <= 32'h00F71E63;
    mem['h0143] <= 32'hFEE44703;
    mem['h0144] <= 32'h01D00793;
    mem['h0145] <= 32'h00E7F863;
    mem['h0146] <= 32'hFEE44703;
    mem['h0147] <= 32'h02000793;
    mem['h0148] <= 32'h04E7F663;
    mem['h0149] <= 32'hFEE44703;
    mem['h014A] <= 32'h01F00793;
    mem['h014B] <= 32'h02F71263;
    mem['h014C] <= 32'hFED44783;
    mem['h014D] <= 32'h00178713;
    mem['h014E] <= 32'hFEF44783;
    mem['h014F] <= 32'h00F75A63;
    mem['h0150] <= 32'hFEF44703;
    mem['h0151] <= 32'hFED44783;
    mem['h0152] <= 32'h00478793;
    mem['h0153] <= 32'h02E7D063;
    mem['h0154] <= 32'hFEE44703;
    mem['h0155] <= 32'h02000793;
    mem['h0156] <= 32'h04F71463;
    mem['h0157] <= 32'hFEF44703;
    mem['h0158] <= 32'hFED44783;
    mem['h0159] <= 32'h00178793;
    mem['h015A] <= 32'h02F71C63;
    mem['h015B] <= 32'hFEF44703;
    mem['h015C] <= 32'h00070793;
    mem['h015D] <= 32'h00279793;
    mem['h015E] <= 32'h00E787B3;
    mem['h015F] <= 32'h00379793;
    mem['h0160] <= 32'h00078713;
    mem['h0161] <= 32'hFEE44783;
    mem['h0162] <= 32'h00F707B3;
    mem['h0163] <= 32'h00279713;
    mem['h0164] <= 32'h052007B7;
    mem['h0165] <= 32'h00F707B3;
    mem['h0166] <= 32'h00200713;
    mem['h0167] <= 32'h00E7A023;
    mem['h0168] <= 32'hFEE44783;
    mem['h0169] <= 32'h00178793;
    mem['h016A] <= 32'hFEF40723;
    mem['h016B] <= 32'hFEE44703;
    mem['h016C] <= 32'h02700793;
    mem['h016D] <= 32'hB6E7FAE3;
    mem['h016E] <= 32'hFEF44783;
    mem['h016F] <= 32'h00178793;
    mem['h0170] <= 32'hFEF407A3;
    mem['h0171] <= 32'hFEF44703;
    mem['h0172] <= 32'h01D00793;
    mem['h0173] <= 32'hB4E7FAE3;
    mem['h0174] <= 32'h00000013;
    mem['h0175] <= 32'h00000013;
    mem['h0176] <= 32'h01C12403;
    mem['h0177] <= 32'h02010113;
    mem['h0178] <= 32'h00008067;
    mem['h0179] <= 32'hFE010113;
    mem['h017A] <= 32'h00812E23;
    mem['h017B] <= 32'h02010413;
    mem['h017C] <= 32'h00B00793;
    mem['h017D] <= 32'hFEF406A3;
    mem['h017E] <= 32'h00300793;
    mem['h017F] <= 32'hFEF40623;
    mem['h0180] <= 32'h02400793;
    mem['h0181] <= 32'hFEF405A3;
    mem['h0182] <= 32'h00E00793;
    mem['h0183] <= 32'hFEF40523;
    mem['h0184] <= 32'hFE0407A3;
    mem['h0185] <= 32'h2010006F;
    mem['h0186] <= 32'hFE040723;
    mem['h0187] <= 32'h1E10006F;
    mem['h0188] <= 32'hFEF44703;
    mem['h0189] <= 32'hFED44783;
    mem['h018A] <= 32'h04F71863;
    mem['h018B] <= 32'hFEE44703;
    mem['h018C] <= 32'hFEC44783;
    mem['h018D] <= 32'h04F76263;
    mem['h018E] <= 32'hFEE44703;
    mem['h018F] <= 32'hFEB44783;
    mem['h0190] <= 32'h02E7EC63;
    mem['h0191] <= 32'hFEF44703;
    mem['h0192] <= 32'h00070793;
    mem['h0193] <= 32'h00279793;
    mem['h0194] <= 32'h00E787B3;
    mem['h0195] <= 32'h00379793;
    mem['h0196] <= 32'h00078713;
    mem['h0197] <= 32'hFEE44783;
    mem['h0198] <= 32'h00F707B3;
    mem['h0199] <= 32'h00279713;
    mem['h019A] <= 32'h052007B7;
    mem['h019B] <= 32'h00F707B3;
    mem['h019C] <= 32'h00A00713;
    mem['h019D] <= 32'h00E7A023;
    mem['h019E] <= 32'hFEE44703;
    mem['h019F] <= 32'h00400793;
    mem['h01A0] <= 32'h04F71A63;
    mem['h01A1] <= 32'hFEF44703;
    mem['h01A2] <= 32'hFEA44783;
    mem['h01A3] <= 32'h04F76463;
    mem['h01A4] <= 32'hFEF44703;
    mem['h01A5] <= 32'hFEA44783;
    mem['h01A6] <= 32'h00478793;
    mem['h01A7] <= 32'h02E7CC63;
    mem['h01A8] <= 32'hFEF44703;
    mem['h01A9] <= 32'h00070793;
    mem['h01AA] <= 32'h00279793;
    mem['h01AB] <= 32'h00E787B3;
    mem['h01AC] <= 32'h00379793;
    mem['h01AD] <= 32'h00078713;
    mem['h01AE] <= 32'hFEE44783;
    mem['h01AF] <= 32'h00F707B3;
    mem['h01B0] <= 32'h00279713;
    mem['h01B1] <= 32'h052007B7;
    mem['h01B2] <= 32'h00F707B3;
    mem['h01B3] <= 32'h00700713;
    mem['h01B4] <= 32'h00E7A023;
    mem['h01B5] <= 32'hFEF44703;
    mem['h01B6] <= 32'hFEA44783;
    mem['h01B7] <= 32'h04F71863;
    mem['h01B8] <= 32'hFEE44703;
    mem['h01B9] <= 32'h00500793;
    mem['h01BA] <= 32'h00F70863;
    mem['h01BB] <= 32'hFEE44703;
    mem['h01BC] <= 32'h00600793;
    mem['h01BD] <= 32'h02F71C63;
    mem['h01BE] <= 32'hFEF44703;
    mem['h01BF] <= 32'h00070793;
    mem['h01C0] <= 32'h00279793;
    mem['h01C1] <= 32'h00E787B3;
    mem['h01C2] <= 32'h00379793;
    mem['h01C3] <= 32'h00078713;
    mem['h01C4] <= 32'hFEE44783;
    mem['h01C5] <= 32'h00F707B3;
    mem['h01C6] <= 32'h00279713;
    mem['h01C7] <= 32'h052007B7;
    mem['h01C8] <= 32'h00F707B3;
    mem['h01C9] <= 32'h00700713;
    mem['h01CA] <= 32'h00E7A023;
    mem['h01CB] <= 32'hFEF44703;
    mem['h01CC] <= 32'hFEA44783;
    mem['h01CD] <= 32'h00478793;
    mem['h01CE] <= 32'h04F71863;
    mem['h01CF] <= 32'hFEE44703;
    mem['h01D0] <= 32'h00500793;
    mem['h01D1] <= 32'h00F70863;
    mem['h01D2] <= 32'hFEE44703;
    mem['h01D3] <= 32'h00600793;
    mem['h01D4] <= 32'h02F71C63;
    mem['h01D5] <= 32'hFEF44703;
    mem['h01D6] <= 32'h00070793;
    mem['h01D7] <= 32'h00279793;
    mem['h01D8] <= 32'h00E787B3;
    mem['h01D9] <= 32'h00379793;
    mem['h01DA] <= 32'h00078713;
    mem['h01DB] <= 32'hFEE44783;
    mem['h01DC] <= 32'h00F707B3;
    mem['h01DD] <= 32'h00279713;
    mem['h01DE] <= 32'h052007B7;
    mem['h01DF] <= 32'h00F707B3;
    mem['h01E0] <= 32'h00700713;
    mem['h01E1] <= 32'h00E7A023;
    mem['h01E2] <= 32'hFEE44703;
    mem['h01E3] <= 32'h00800793;
    mem['h01E4] <= 32'h04F71A63;
    mem['h01E5] <= 32'hFEF44703;
    mem['h01E6] <= 32'hFEA44783;
    mem['h01E7] <= 32'h04F76463;
    mem['h01E8] <= 32'hFEF44703;
    mem['h01E9] <= 32'hFEA44783;
    mem['h01EA] <= 32'h00478793;
    mem['h01EB] <= 32'h02E7CC63;
    mem['h01EC] <= 32'hFEF44703;
    mem['h01ED] <= 32'h00070793;
    mem['h01EE] <= 32'h00279793;
    mem['h01EF] <= 32'h00E787B3;
    mem['h01F0] <= 32'h00379793;
    mem['h01F1] <= 32'h00078713;
    mem['h01F2] <= 32'hFEE44783;
    mem['h01F3] <= 32'h00F707B3;
    mem['h01F4] <= 32'h00279713;
    mem['h01F5] <= 32'h052007B7;
    mem['h01F6] <= 32'h00F707B3;
    mem['h01F7] <= 32'h00700713;
    mem['h01F8] <= 32'h00E7A023;
    mem['h01F9] <= 32'hFEF44703;
    mem['h01FA] <= 32'hFEA44783;
    mem['h01FB] <= 32'h00278793;
    mem['h01FC] <= 32'h04F71863;
    mem['h01FD] <= 32'hFEE44703;
    mem['h01FE] <= 32'h00900793;
    mem['h01FF] <= 32'h00F70863;
    mem['h0200] <= 32'hFEE44703;
    mem['h0201] <= 32'h00A00793;
    mem['h0202] <= 32'h02F71C63;
    mem['h0203] <= 32'hFEF44703;
    mem['h0204] <= 32'h00070793;
    mem['h0205] <= 32'h00279793;
    mem['h0206] <= 32'h00E787B3;
    mem['h0207] <= 32'h00379793;
    mem['h0208] <= 32'h00078713;
    mem['h0209] <= 32'hFEE44783;
    mem['h020A] <= 32'h00F707B3;
    mem['h020B] <= 32'h00279713;
    mem['h020C] <= 32'h052007B7;
    mem['h020D] <= 32'h00F707B3;
    mem['h020E] <= 32'h00700713;
    mem['h020F] <= 32'h00E7A023;
    mem['h0210] <= 32'hFEE44703;
    mem['h0211] <= 32'h00A00793;
    mem['h0212] <= 32'h04F71C63;
    mem['h0213] <= 32'hFEA44783;
    mem['h0214] <= 32'h00178713;
    mem['h0215] <= 32'hFEF44783;
    mem['h0216] <= 32'h04F75463;
    mem['h0217] <= 32'hFEF44703;
    mem['h0218] <= 32'hFEA44783;
    mem['h0219] <= 32'h00478793;
    mem['h021A] <= 32'h02E7CC63;
    mem['h021B] <= 32'hFEF44703;
    mem['h021C] <= 32'h00070793;
    mem['h021D] <= 32'h00279793;
    mem['h021E] <= 32'h00E787B3;
    mem['h021F] <= 32'h00379793;
    mem['h0220] <= 32'h00078713;
    mem['h0221] <= 32'hFEE44783;
    mem['h0222] <= 32'h00F707B3;
    mem['h0223] <= 32'h00279713;
    mem['h0224] <= 32'h052007B7;
    mem['h0225] <= 32'h00F707B3;
    mem['h0226] <= 32'h00700713;
    mem['h0227] <= 32'h00E7A023;
    mem['h0228] <= 32'hFEE44703;
    mem['h0229] <= 32'h00C00793;
    mem['h022A] <= 32'h04F71C63;
    mem['h022B] <= 32'hFEA44783;
    mem['h022C] <= 32'h00178713;
    mem['h022D] <= 32'hFEF44783;
    mem['h022E] <= 32'h04F75463;
    mem['h022F] <= 32'hFEF44703;
    mem['h0230] <= 32'hFEA44783;
    mem['h0231] <= 32'h00478793;
    mem['h0232] <= 32'h02E7CC63;
    mem['h0233] <= 32'hFEF44703;
    mem['h0234] <= 32'h00070793;
    mem['h0235] <= 32'h00279793;
    mem['h0236] <= 32'h00E787B3;
    mem['h0237] <= 32'h00379793;
    mem['h0238] <= 32'h00078713;
    mem['h0239] <= 32'hFEE44783;
    mem['h023A] <= 32'h00F707B3;
    mem['h023B] <= 32'h00279713;
    mem['h023C] <= 32'h052007B7;
    mem['h023D] <= 32'h00F707B3;
    mem['h023E] <= 32'h00700713;
    mem['h023F] <= 32'h00E7A023;
    mem['h0240] <= 32'hFEE44703;
    mem['h0241] <= 32'h00C00793;
    mem['h0242] <= 32'h04F71263;
    mem['h0243] <= 32'hFEF44703;
    mem['h0244] <= 32'hFEA44783;
    mem['h0245] <= 32'h02F71C63;
    mem['h0246] <= 32'hFEF44703;
    mem['h0247] <= 32'h00070793;
    mem['h0248] <= 32'h00279793;
    mem['h0249] <= 32'h00E787B3;
    mem['h024A] <= 32'h00379793;
    mem['h024B] <= 32'h00078713;
    mem['h024C] <= 32'hFEE44783;
    mem['h024D] <= 32'h00F707B3;
    mem['h024E] <= 32'h00279713;
    mem['h024F] <= 32'h052007B7;
    mem['h0250] <= 32'h00F707B3;
    mem['h0251] <= 32'h00700713;
    mem['h0252] <= 32'h00E7A023;
    mem['h0253] <= 32'hFEE44703;
    mem['h0254] <= 32'h00E00793;
    mem['h0255] <= 32'h04F71A63;
    mem['h0256] <= 32'hFEF44703;
    mem['h0257] <= 32'hFEA44783;
    mem['h0258] <= 32'h04F76463;
    mem['h0259] <= 32'hFEF44703;
    mem['h025A] <= 32'hFEA44783;
    mem['h025B] <= 32'h00478793;
    mem['h025C] <= 32'h02E7CC63;
    mem['h025D] <= 32'hFEF44703;
    mem['h025E] <= 32'h00070793;
    mem['h025F] <= 32'h00279793;
    mem['h0260] <= 32'h00E787B3;
    mem['h0261] <= 32'h00379793;
    mem['h0262] <= 32'h00078713;
    mem['h0263] <= 32'hFEE44783;
    mem['h0264] <= 32'h00F707B3;
    mem['h0265] <= 32'h00279713;
    mem['h0266] <= 32'h052007B7;
    mem['h0267] <= 32'h00F707B3;
    mem['h0268] <= 32'h00700713;
    mem['h0269] <= 32'h00E7A023;
    mem['h026A] <= 32'hFEE44703;
    mem['h026B] <= 32'h01000793;
    mem['h026C] <= 32'h04F71C63;
    mem['h026D] <= 32'hFEA44783;
    mem['h026E] <= 32'h00178713;
    mem['h026F] <= 32'hFEF44783;
    mem['h0270] <= 32'h04F75463;
    mem['h0271] <= 32'hFEF44703;
    mem['h0272] <= 32'hFEA44783;
    mem['h0273] <= 32'h00478793;
    mem['h0274] <= 32'h02E7CC63;
    mem['h0275] <= 32'hFEF44703;
    mem['h0276] <= 32'h00070793;
    mem['h0277] <= 32'h00279793;
    mem['h0278] <= 32'h00E787B3;
    mem['h0279] <= 32'h00379793;
    mem['h027A] <= 32'h00078713;
    mem['h027B] <= 32'hFEE44783;
    mem['h027C] <= 32'h00F707B3;
    mem['h027D] <= 32'h00279713;
    mem['h027E] <= 32'h052007B7;
    mem['h027F] <= 32'h00F707B3;
    mem['h0280] <= 32'h00700713;
    mem['h0281] <= 32'h00E7A023;
    mem['h0282] <= 32'hFEE44703;
    mem['h0283] <= 32'h01000793;
    mem['h0284] <= 32'h04F71263;
    mem['h0285] <= 32'hFEF44703;
    mem['h0286] <= 32'hFEA44783;
    mem['h0287] <= 32'h02F71C63;
    mem['h0288] <= 32'hFEF44703;
    mem['h0289] <= 32'h00070793;
    mem['h028A] <= 32'h00279793;
    mem['h028B] <= 32'h00E787B3;
    mem['h028C] <= 32'h00379793;
    mem['h028D] <= 32'h00078713;
    mem['h028E] <= 32'hFEE44783;
    mem['h028F] <= 32'h00F707B3;
    mem['h0290] <= 32'h00279713;
    mem['h0291] <= 32'h052007B7;
    mem['h0292] <= 32'h00F707B3;
    mem['h0293] <= 32'h00700713;
    mem['h0294] <= 32'h00E7A023;
    mem['h0295] <= 32'hFEE44703;
    mem['h0296] <= 32'h01300793;
    mem['h0297] <= 32'h04F71A63;
    mem['h0298] <= 32'hFEF44703;
    mem['h0299] <= 32'hFEA44783;
    mem['h029A] <= 32'h04F76463;
    mem['h029B] <= 32'hFEF44703;
    mem['h029C] <= 32'hFEA44783;
    mem['h029D] <= 32'h00478793;
    mem['h029E] <= 32'h02E7CC63;
    mem['h029F] <= 32'hFEF44703;
    mem['h02A0] <= 32'h00070793;
    mem['h02A1] <= 32'h00279793;
    mem['h02A2] <= 32'h00E787B3;
    mem['h02A3] <= 32'h00379793;
    mem['h02A4] <= 32'h00078713;
    mem['h02A5] <= 32'hFEE44783;
    mem['h02A6] <= 32'h00F707B3;
    mem['h02A7] <= 32'h00279713;
    mem['h02A8] <= 32'h052007B7;
    mem['h02A9] <= 32'h00F707B3;
    mem['h02AA] <= 32'h00A00713;
    mem['h02AB] <= 32'h00E7A023;
    mem['h02AC] <= 32'hFEF44703;
    mem['h02AD] <= 32'hFEA44783;
    mem['h02AE] <= 32'h04F71863;
    mem['h02AF] <= 32'hFEE44703;
    mem['h02B0] <= 32'h01400793;
    mem['h02B1] <= 32'h00F70863;
    mem['h02B2] <= 32'hFEE44703;
    mem['h02B3] <= 32'h01500793;
    mem['h02B4] <= 32'h02F71C63;
    mem['h02B5] <= 32'hFEF44703;
    mem['h02B6] <= 32'h00070793;
    mem['h02B7] <= 32'h00279793;
    mem['h02B8] <= 32'h00E787B3;
    mem['h02B9] <= 32'h00379793;
    mem['h02BA] <= 32'h00078713;
    mem['h02BB] <= 32'hFEE44783;
    mem['h02BC] <= 32'h00F707B3;
    mem['h02BD] <= 32'h00279713;
    mem['h02BE] <= 32'h052007B7;
    mem['h02BF] <= 32'h00F707B3;
    mem['h02C0] <= 32'h00A00713;
    mem['h02C1] <= 32'h00E7A023;
    mem['h02C2] <= 32'hFEF44703;
    mem['h02C3] <= 32'hFEA44783;
    mem['h02C4] <= 32'h00478793;
    mem['h02C5] <= 32'h04F71863;
    mem['h02C6] <= 32'hFEE44703;
    mem['h02C7] <= 32'h01400793;
    mem['h02C8] <= 32'h00F70863;
    mem['h02C9] <= 32'hFEE44703;
    mem['h02CA] <= 32'h01500793;
    mem['h02CB] <= 32'h02F71C63;
    mem['h02CC] <= 32'hFEF44703;
    mem['h02CD] <= 32'h00070793;
    mem['h02CE] <= 32'h00279793;
    mem['h02CF] <= 32'h00E787B3;
    mem['h02D0] <= 32'h00379793;
    mem['h02D1] <= 32'h00078713;
    mem['h02D2] <= 32'hFEE44783;
    mem['h02D3] <= 32'h00F707B3;
    mem['h02D4] <= 32'h00279713;
    mem['h02D5] <= 32'h052007B7;
    mem['h02D6] <= 32'h00F707B3;
    mem['h02D7] <= 32'h00A00713;
    mem['h02D8] <= 32'h00E7A023;
    mem['h02D9] <= 32'hFEE44703;
    mem['h02DA] <= 32'h01700793;
    mem['h02DB] <= 32'h04F71A63;
    mem['h02DC] <= 32'hFEF44703;
    mem['h02DD] <= 32'hFEA44783;
    mem['h02DE] <= 32'h04F76463;
    mem['h02DF] <= 32'hFEF44703;
    mem['h02E0] <= 32'hFEA44783;
    mem['h02E1] <= 32'h00478793;
    mem['h02E2] <= 32'h02E7CC63;
    mem['h02E3] <= 32'hFEF44703;
    mem['h02E4] <= 32'h00070793;
    mem['h02E5] <= 32'h00279793;
    mem['h02E6] <= 32'h00E787B3;
    mem['h02E7] <= 32'h00379793;
    mem['h02E8] <= 32'h00078713;
    mem['h02E9] <= 32'hFEE44783;
    mem['h02EA] <= 32'h00F707B3;
    mem['h02EB] <= 32'h00279713;
    mem['h02EC] <= 32'h052007B7;
    mem['h02ED] <= 32'h00F707B3;
    mem['h02EE] <= 32'h00A00713;
    mem['h02EF] <= 32'h00E7A023;
    mem['h02F0] <= 32'hFEF44703;
    mem['h02F1] <= 32'hFEA44783;
    mem['h02F2] <= 32'h00278793;
    mem['h02F3] <= 32'h04F71863;
    mem['h02F4] <= 32'hFEE44703;
    mem['h02F5] <= 32'h01800793;
    mem['h02F6] <= 32'h00F70863;
    mem['h02F7] <= 32'hFEE44703;
    mem['h02F8] <= 32'h01900793;
    mem['h02F9] <= 32'h02F71C63;
    mem['h02FA] <= 32'hFEF44703;
    mem['h02FB] <= 32'h00070793;
    mem['h02FC] <= 32'h00279793;
    mem['h02FD] <= 32'h00E787B3;
    mem['h02FE] <= 32'h00379793;
    mem['h02FF] <= 32'h00078713;
    mem['h0300] <= 32'hFEE44783;
    mem['h0301] <= 32'h00F707B3;
    mem['h0302] <= 32'h00279713;
    mem['h0303] <= 32'h052007B7;
    mem['h0304] <= 32'h00F707B3;
    mem['h0305] <= 32'h00A00713;
    mem['h0306] <= 32'h00E7A023;
    mem['h0307] <= 32'hFEE44703;
    mem['h0308] <= 32'h01900793;
    mem['h0309] <= 32'h04F71A63;
    mem['h030A] <= 32'hFEF44703;
    mem['h030B] <= 32'hFEA44783;
    mem['h030C] <= 32'h04F76463;
    mem['h030D] <= 32'hFEF44703;
    mem['h030E] <= 32'hFEA44783;
    mem['h030F] <= 32'h00478793;
    mem['h0310] <= 32'h02E7CC63;
    mem['h0311] <= 32'hFEF44703;
    mem['h0312] <= 32'h00070793;
    mem['h0313] <= 32'h00279793;
    mem['h0314] <= 32'h00E787B3;
    mem['h0315] <= 32'h00379793;
    mem['h0316] <= 32'h00078713;
    mem['h0317] <= 32'hFEE44783;
    mem['h0318] <= 32'h00F707B3;
    mem['h0319] <= 32'h00279713;
    mem['h031A] <= 32'h052007B7;
    mem['h031B] <= 32'h00F707B3;
    mem['h031C] <= 32'h00A00713;
    mem['h031D] <= 32'h00E7A023;
    mem['h031E] <= 32'hFEE44703;
    mem['h031F] <= 32'h01B00793;
    mem['h0320] <= 32'h04F71A63;
    mem['h0321] <= 32'hFEF44703;
    mem['h0322] <= 32'hFEA44783;
    mem['h0323] <= 32'h04F76463;
    mem['h0324] <= 32'hFEF44703;
    mem['h0325] <= 32'hFEA44783;
    mem['h0326] <= 32'h00478793;
    mem['h0327] <= 32'h02E7CC63;
    mem['h0328] <= 32'hFEF44703;
    mem['h0329] <= 32'h00070793;
    mem['h032A] <= 32'h00279793;
    mem['h032B] <= 32'h00E787B3;
    mem['h032C] <= 32'h00379793;
    mem['h032D] <= 32'h00078713;
    mem['h032E] <= 32'hFEE44783;
    mem['h032F] <= 32'h00F707B3;
    mem['h0330] <= 32'h00279713;
    mem['h0331] <= 32'h052007B7;
    mem['h0332] <= 32'h00F707B3;
    mem['h0333] <= 32'h00A00713;
    mem['h0334] <= 32'h00E7A023;
    mem['h0335] <= 32'hFEE44703;
    mem['h0336] <= 32'h01D00793;
    mem['h0337] <= 32'h04F71A63;
    mem['h0338] <= 32'hFEF44703;
    mem['h0339] <= 32'hFEA44783;
    mem['h033A] <= 32'h04F76463;
    mem['h033B] <= 32'hFEF44703;
    mem['h033C] <= 32'hFEA44783;
    mem['h033D] <= 32'h00478793;
    mem['h033E] <= 32'h02E7CC63;
    mem['h033F] <= 32'hFEF44703;
    mem['h0340] <= 32'h00070793;
    mem['h0341] <= 32'h00279793;
    mem['h0342] <= 32'h00E787B3;
    mem['h0343] <= 32'h00379793;
    mem['h0344] <= 32'h00078713;
    mem['h0345] <= 32'hFEE44783;
    mem['h0346] <= 32'h00F707B3;
    mem['h0347] <= 32'h00279713;
    mem['h0348] <= 32'h052007B7;
    mem['h0349] <= 32'h00F707B3;
    mem['h034A] <= 32'h00A00713;
    mem['h034B] <= 32'h00E7A023;
    mem['h034C] <= 32'hFEF44703;
    mem['h034D] <= 32'hFEA44783;
    mem['h034E] <= 32'h04F71863;
    mem['h034F] <= 32'hFEE44703;
    mem['h0350] <= 32'h01E00793;
    mem['h0351] <= 32'h00F70863;
    mem['h0352] <= 32'hFEE44703;
    mem['h0353] <= 32'h01F00793;
    mem['h0354] <= 32'h02F71C63;
    mem['h0355] <= 32'hFEF44703;
    mem['h0356] <= 32'h00070793;
    mem['h0357] <= 32'h00279793;
    mem['h0358] <= 32'h00E787B3;
    mem['h0359] <= 32'h00379793;
    mem['h035A] <= 32'h00078713;
    mem['h035B] <= 32'hFEE44783;
    mem['h035C] <= 32'h00F707B3;
    mem['h035D] <= 32'h00279713;
    mem['h035E] <= 32'h052007B7;
    mem['h035F] <= 32'h00F707B3;
    mem['h0360] <= 32'h00A00713;
    mem['h0361] <= 32'h00E7A023;
    mem['h0362] <= 32'hFEF44703;
    mem['h0363] <= 32'hFEA44783;
    mem['h0364] <= 32'h00278793;
    mem['h0365] <= 32'h04F71863;
    mem['h0366] <= 32'hFEE44703;
    mem['h0367] <= 32'h01E00793;
    mem['h0368] <= 32'h00F70863;
    mem['h0369] <= 32'hFEE44703;
    mem['h036A] <= 32'h01F00793;
    mem['h036B] <= 32'h02F71C63;
    mem['h036C] <= 32'hFEF44703;
    mem['h036D] <= 32'h00070793;
    mem['h036E] <= 32'h00279793;
    mem['h036F] <= 32'h00E787B3;
    mem['h0370] <= 32'h00379793;
    mem['h0371] <= 32'h00078713;
    mem['h0372] <= 32'hFEE44783;
    mem['h0373] <= 32'h00F707B3;
    mem['h0374] <= 32'h00279713;
    mem['h0375] <= 32'h052007B7;
    mem['h0376] <= 32'h00F707B3;
    mem['h0377] <= 32'h00A00713;
    mem['h0378] <= 32'h00E7A023;
    mem['h0379] <= 32'hFEE44703;
    mem['h037A] <= 32'h01F00793;
    mem['h037B] <= 32'h04F71A63;
    mem['h037C] <= 32'hFEF44703;
    mem['h037D] <= 32'hFEA44783;
    mem['h037E] <= 32'h04F76463;
    mem['h037F] <= 32'hFEF44703;
    mem['h0380] <= 32'hFEA44783;
    mem['h0381] <= 32'h00278793;
    mem['h0382] <= 32'h02E7CC63;
    mem['h0383] <= 32'hFEF44703;
    mem['h0384] <= 32'h00070793;
    mem['h0385] <= 32'h00279793;
    mem['h0386] <= 32'h00E787B3;
    mem['h0387] <= 32'h00379793;
    mem['h0388] <= 32'h00078713;
    mem['h0389] <= 32'hFEE44783;
    mem['h038A] <= 32'h00F707B3;
    mem['h038B] <= 32'h00279713;
    mem['h038C] <= 32'h052007B7;
    mem['h038D] <= 32'h00F707B3;
    mem['h038E] <= 32'h00A00713;
    mem['h038F] <= 32'h00E7A023;
    mem['h0390] <= 32'hFEF44703;
    mem['h0391] <= 32'hFEA44783;
    mem['h0392] <= 32'h04F71863;
    mem['h0393] <= 32'hFEE44703;
    mem['h0394] <= 32'h02000793;
    mem['h0395] <= 32'h04E7F263;
    mem['h0396] <= 32'hFEE44703;
    mem['h0397] <= 32'h02300793;
    mem['h0398] <= 32'h02E7EC63;
    mem['h0399] <= 32'hFEF44703;
    mem['h039A] <= 32'h00070793;
    mem['h039B] <= 32'h00279793;
    mem['h039C] <= 32'h00E787B3;
    mem['h039D] <= 32'h00379793;
    mem['h039E] <= 32'h00078713;
    mem['h039F] <= 32'hFEE44783;
    mem['h03A0] <= 32'h00F707B3;
    mem['h03A1] <= 32'h00279713;
    mem['h03A2] <= 32'h052007B7;
    mem['h03A3] <= 32'h00F707B3;
    mem['h03A4] <= 32'h00A00713;
    mem['h03A5] <= 32'h00E7A023;
    mem['h03A6] <= 32'hFEF44703;
    mem['h03A7] <= 32'hFEA44783;
    mem['h03A8] <= 32'h00278793;
    mem['h03A9] <= 32'h04F71863;
    mem['h03AA] <= 32'hFEE44703;
    mem['h03AB] <= 32'h02000793;
    mem['h03AC] <= 32'h04E7F263;
    mem['h03AD] <= 32'hFEE44703;
    mem['h03AE] <= 32'h02300793;
    mem['h03AF] <= 32'h02E7EC63;
    mem['h03B0] <= 32'hFEF44703;
    mem['h03B1] <= 32'h00070793;
    mem['h03B2] <= 32'h00279793;
    mem['h03B3] <= 32'h00E787B3;
    mem['h03B4] <= 32'h00379793;
    mem['h03B5] <= 32'h00078713;
    mem['h03B6] <= 32'hFEE44783;
    mem['h03B7] <= 32'h00F707B3;
    mem['h03B8] <= 32'h00279713;
    mem['h03B9] <= 32'h052007B7;
    mem['h03BA] <= 32'h00F707B3;
    mem['h03BB] <= 32'h00A00713;
    mem['h03BC] <= 32'h00E7A023;
    mem['h03BD] <= 32'hFEF44703;
    mem['h03BE] <= 32'hFEA44783;
    mem['h03BF] <= 32'h00478793;
    mem['h03C0] <= 32'h04F71863;
    mem['h03C1] <= 32'hFEE44703;
    mem['h03C2] <= 32'h02000793;
    mem['h03C3] <= 32'h04E7F263;
    mem['h03C4] <= 32'hFEE44703;
    mem['h03C5] <= 32'h02300793;
    mem['h03C6] <= 32'h02E7EC63;
    mem['h03C7] <= 32'hFEF44703;
    mem['h03C8] <= 32'h00070793;
    mem['h03C9] <= 32'h00279793;
    mem['h03CA] <= 32'h00E787B3;
    mem['h03CB] <= 32'h00379793;
    mem['h03CC] <= 32'h00078713;
    mem['h03CD] <= 32'hFEE44783;
    mem['h03CE] <= 32'h00F707B3;
    mem['h03CF] <= 32'h00279713;
    mem['h03D0] <= 32'h052007B7;
    mem['h03D1] <= 32'h00F707B3;
    mem['h03D2] <= 32'h00A00713;
    mem['h03D3] <= 32'h00E7A023;
    mem['h03D4] <= 32'hFEE44703;
    mem['h03D5] <= 32'h02100793;
    mem['h03D6] <= 32'h04F71463;
    mem['h03D7] <= 32'hFEF44703;
    mem['h03D8] <= 32'hFEA44783;
    mem['h03D9] <= 32'h00178793;
    mem['h03DA] <= 32'h02F71C63;
    mem['h03DB] <= 32'hFEF44703;
    mem['h03DC] <= 32'h00070793;
    mem['h03DD] <= 32'h00279793;
    mem['h03DE] <= 32'h00E787B3;
    mem['h03DF] <= 32'h00379793;
    mem['h03E0] <= 32'h00078713;
    mem['h03E1] <= 32'hFEE44783;
    mem['h03E2] <= 32'h00F707B3;
    mem['h03E3] <= 32'h00279713;
    mem['h03E4] <= 32'h052007B7;
    mem['h03E5] <= 32'h00F707B3;
    mem['h03E6] <= 32'h00A00713;
    mem['h03E7] <= 32'h00E7A023;
    mem['h03E8] <= 32'hFEE44703;
    mem['h03E9] <= 32'h02300793;
    mem['h03EA] <= 32'h04F71463;
    mem['h03EB] <= 32'hFEF44703;
    mem['h03EC] <= 32'hFEA44783;
    mem['h03ED] <= 32'h00378793;
    mem['h03EE] <= 32'h02F71C63;
    mem['h03EF] <= 32'hFEF44703;
    mem['h03F0] <= 32'h00070793;
    mem['h03F1] <= 32'h00279793;
    mem['h03F2] <= 32'h00E787B3;
    mem['h03F3] <= 32'h00379793;
    mem['h03F4] <= 32'h00078713;
    mem['h03F5] <= 32'hFEE44783;
    mem['h03F6] <= 32'h00F707B3;
    mem['h03F7] <= 32'h00279713;
    mem['h03F8] <= 32'h052007B7;
    mem['h03F9] <= 32'h00F707B3;
    mem['h03FA] <= 32'h00A00713;
    mem['h03FB] <= 32'h00E7A023;
    mem['h03FC] <= 32'hFEE44783;
    mem['h03FD] <= 32'h00178793;
    mem['h03FE] <= 32'hFEF40723;
    mem['h03FF] <= 32'hFEE44703;
    mem['h0400] <= 32'h02700793;
    mem['h0401] <= 32'hE0E7FE63;
    mem['h0402] <= 32'hFEF44783;
    mem['h0403] <= 32'h00178793;
    mem['h0404] <= 32'hFEF407A3;
    mem['h0405] <= 32'hFEF44703;
    mem['h0406] <= 32'h01D00793;
    mem['h0407] <= 32'hDEE7FE63;
    mem['h0408] <= 32'h00000013;
    mem['h0409] <= 32'h00000013;
    mem['h040A] <= 32'h01C12403;
    mem['h040B] <= 32'h02010113;
    mem['h040C] <= 32'h00008067;
    mem['h040D] <= 32'hFE010113;
    mem['h040E] <= 32'h00812E23;
    mem['h040F] <= 32'h02010413;
    mem['h0410] <= 32'h01600793;
    mem['h0411] <= 32'hFEF406A3;
    mem['h0412] <= 32'hFE0407A3;
    mem['h0413] <= 32'h2450006F;
    mem['h0414] <= 32'hFE040723;
    mem['h0415] <= 32'h2250006F;
    mem['h0416] <= 32'hFEF44703;
    mem['h0417] <= 32'hFED44783;
    mem['h0418] <= 32'h04F71863;
    mem['h0419] <= 32'hFEE44703;
    mem['h041A] <= 32'h00200793;
    mem['h041B] <= 32'h04E7F263;
    mem['h041C] <= 32'hFEE44703;
    mem['h041D] <= 32'h00500793;
    mem['h041E] <= 32'h02E7EC63;
    mem['h041F] <= 32'hFEF44703;
    mem['h0420] <= 32'h00070793;
    mem['h0421] <= 32'h00279793;
    mem['h0422] <= 32'h00E787B3;
    mem['h0423] <= 32'h00379793;
    mem['h0424] <= 32'h00078713;
    mem['h0425] <= 32'hFEE44783;
    mem['h0426] <= 32'h00F707B3;
    mem['h0427] <= 32'h00279713;
    mem['h0428] <= 32'h052007B7;
    mem['h0429] <= 32'h00F707B3;
    mem['h042A] <= 32'h00200713;
    mem['h042B] <= 32'h00E7A023;
    mem['h042C] <= 32'hFEE44703;
    mem['h042D] <= 32'h00400793;
    mem['h042E] <= 32'h04F71A63;
    mem['h042F] <= 32'hFEF44703;
    mem['h0430] <= 32'hFED44783;
    mem['h0431] <= 32'h04F76463;
    mem['h0432] <= 32'hFEF44703;
    mem['h0433] <= 32'hFED44783;
    mem['h0434] <= 32'h00478793;
    mem['h0435] <= 32'h02E7CC63;
    mem['h0436] <= 32'hFEF44703;
    mem['h0437] <= 32'h00070793;
    mem['h0438] <= 32'h00279793;
    mem['h0439] <= 32'h00E787B3;
    mem['h043A] <= 32'h00379793;
    mem['h043B] <= 32'h00078713;
    mem['h043C] <= 32'hFEE44783;
    mem['h043D] <= 32'h00F707B3;
    mem['h043E] <= 32'h00279713;
    mem['h043F] <= 32'h052007B7;
    mem['h0440] <= 32'h00F707B3;
    mem['h0441] <= 32'h00200713;
    mem['h0442] <= 32'h00E7A023;
    mem['h0443] <= 32'hFEE44703;
    mem['h0444] <= 32'h00700793;
    mem['h0445] <= 32'h04F71A63;
    mem['h0446] <= 32'hFEF44703;
    mem['h0447] <= 32'hFED44783;
    mem['h0448] <= 32'h04F76463;
    mem['h0449] <= 32'hFEF44703;
    mem['h044A] <= 32'hFED44783;
    mem['h044B] <= 32'h00478793;
    mem['h044C] <= 32'h02E7CC63;
    mem['h044D] <= 32'hFEF44703;
    mem['h044E] <= 32'h00070793;
    mem['h044F] <= 32'h00279793;
    mem['h0450] <= 32'h00E787B3;
    mem['h0451] <= 32'h00379793;
    mem['h0452] <= 32'h00078713;
    mem['h0453] <= 32'hFEE44783;
    mem['h0454] <= 32'h00F707B3;
    mem['h0455] <= 32'h00279713;
    mem['h0456] <= 32'h052007B7;
    mem['h0457] <= 32'h00F707B3;
    mem['h0458] <= 32'h00200713;
    mem['h0459] <= 32'h00E7A023;
    mem['h045A] <= 32'hFEE44703;
    mem['h045B] <= 32'h00800793;
    mem['h045C] <= 32'h06F71263;
    mem['h045D] <= 32'hFEF44703;
    mem['h045E] <= 32'hFED44783;
    mem['h045F] <= 32'h02F70263;
    mem['h0460] <= 32'hFEF44703;
    mem['h0461] <= 32'hFED44783;
    mem['h0462] <= 32'h00278793;
    mem['h0463] <= 32'h00F70A63;
    mem['h0464] <= 32'hFEF44703;
    mem['h0465] <= 32'hFED44783;
    mem['h0466] <= 32'h00478793;
    mem['h0467] <= 32'h02F71C63;
    mem['h0468] <= 32'hFEF44703;
    mem['h0469] <= 32'h00070793;
    mem['h046A] <= 32'h00279793;
    mem['h046B] <= 32'h00E787B3;
    mem['h046C] <= 32'h00379793;
    mem['h046D] <= 32'h00078713;
    mem['h046E] <= 32'hFEE44783;
    mem['h046F] <= 32'h00F707B3;
    mem['h0470] <= 32'h00279713;
    mem['h0471] <= 32'h052007B7;
    mem['h0472] <= 32'h00F707B3;
    mem['h0473] <= 32'h00200713;
    mem['h0474] <= 32'h00E7A023;
    mem['h0475] <= 32'hFEF44703;
    mem['h0476] <= 32'hFED44783;
    mem['h0477] <= 32'h04F71863;
    mem['h0478] <= 32'hFEE44703;
    mem['h0479] <= 32'h00900793;
    mem['h047A] <= 32'h04E7F263;
    mem['h047B] <= 32'hFEE44703;
    mem['h047C] <= 32'h00C00793;
    mem['h047D] <= 32'h02E7EC63;
    mem['h047E] <= 32'hFEF44703;
    mem['h047F] <= 32'h00070793;
    mem['h0480] <= 32'h00279793;
    mem['h0481] <= 32'h00E787B3;
    mem['h0482] <= 32'h00379793;
    mem['h0483] <= 32'h00078713;
    mem['h0484] <= 32'hFEE44783;
    mem['h0485] <= 32'h00F707B3;
    mem['h0486] <= 32'h00279713;
    mem['h0487] <= 32'h052007B7;
    mem['h0488] <= 32'h00F707B3;
    mem['h0489] <= 32'h00200713;
    mem['h048A] <= 32'h00E7A023;
    mem['h048B] <= 32'hFEE44703;
    mem['h048C] <= 32'h00B00793;
    mem['h048D] <= 32'h04F71A63;
    mem['h048E] <= 32'hFEF44703;
    mem['h048F] <= 32'hFED44783;
    mem['h0490] <= 32'h04F76463;
    mem['h0491] <= 32'hFEF44703;
    mem['h0492] <= 32'hFED44783;
    mem['h0493] <= 32'h00478793;
    mem['h0494] <= 32'h02E7CC63;
    mem['h0495] <= 32'hFEF44703;
    mem['h0496] <= 32'h00070793;
    mem['h0497] <= 32'h00279793;
    mem['h0498] <= 32'h00E787B3;
    mem['h0499] <= 32'h00379793;
    mem['h049A] <= 32'h00078713;
    mem['h049B] <= 32'hFEE44783;
    mem['h049C] <= 32'h00F707B3;
    mem['h049D] <= 32'h00279713;
    mem['h049E] <= 32'h052007B7;
    mem['h049F] <= 32'h00F707B3;
    mem['h04A0] <= 32'h00200713;
    mem['h04A1] <= 32'h00E7A023;
    mem['h04A2] <= 32'hFEE44703;
    mem['h04A3] <= 32'h00E00793;
    mem['h04A4] <= 32'h04F71A63;
    mem['h04A5] <= 32'hFEF44703;
    mem['h04A6] <= 32'hFED44783;
    mem['h04A7] <= 32'h04F76463;
    mem['h04A8] <= 32'hFEF44703;
    mem['h04A9] <= 32'hFED44783;
    mem['h04AA] <= 32'h00478793;
    mem['h04AB] <= 32'h02E7CC63;
    mem['h04AC] <= 32'hFEF44703;
    mem['h04AD] <= 32'h00070793;
    mem['h04AE] <= 32'h00279793;
    mem['h04AF] <= 32'h00E787B3;
    mem['h04B0] <= 32'h00379793;
    mem['h04B1] <= 32'h00078713;
    mem['h04B2] <= 32'hFEE44783;
    mem['h04B3] <= 32'h00F707B3;
    mem['h04B4] <= 32'h00279713;
    mem['h04B5] <= 32'h052007B7;
    mem['h04B6] <= 32'h00F707B3;
    mem['h04B7] <= 32'h00200713;
    mem['h04B8] <= 32'h00E7A023;
    mem['h04B9] <= 32'hFEE44703;
    mem['h04BA] <= 32'h00F00793;
    mem['h04BB] <= 32'h04F71263;
    mem['h04BC] <= 32'hFEF44703;
    mem['h04BD] <= 32'hFED44783;
    mem['h04BE] <= 32'h02F71C63;
    mem['h04BF] <= 32'hFEF44703;
    mem['h04C0] <= 32'h00070793;
    mem['h04C1] <= 32'h00279793;
    mem['h04C2] <= 32'h00E787B3;
    mem['h04C3] <= 32'h00379793;
    mem['h04C4] <= 32'h00078713;
    mem['h04C5] <= 32'hFEE44783;
    mem['h04C6] <= 32'h00F707B3;
    mem['h04C7] <= 32'h00279713;
    mem['h04C8] <= 32'h052007B7;
    mem['h04C9] <= 32'h00F707B3;
    mem['h04CA] <= 32'h00200713;
    mem['h04CB] <= 32'h00E7A023;
    mem['h04CC] <= 32'hFEE44703;
    mem['h04CD] <= 32'h01000793;
    mem['h04CE] <= 32'h04F71463;
    mem['h04CF] <= 32'hFEF44703;
    mem['h04D0] <= 32'hFED44783;
    mem['h04D1] <= 32'h00178793;
    mem['h04D2] <= 32'h02F71C63;
    mem['h04D3] <= 32'hFEF44703;
    mem['h04D4] <= 32'h00070793;
    mem['h04D5] <= 32'h00279793;
    mem['h04D6] <= 32'h00E787B3;
    mem['h04D7] <= 32'h00379793;
    mem['h04D8] <= 32'h00078713;
    mem['h04D9] <= 32'hFEE44783;
    mem['h04DA] <= 32'h00F707B3;
    mem['h04DB] <= 32'h00279713;
    mem['h04DC] <= 32'h052007B7;
    mem['h04DD] <= 32'h00F707B3;
    mem['h04DE] <= 32'h00200713;
    mem['h04DF] <= 32'h00E7A023;
    mem['h04E0] <= 32'hFEE44703;
    mem['h04E1] <= 32'h00F00793;
    mem['h04E2] <= 32'h04F71463;
    mem['h04E3] <= 32'hFEF44703;
    mem['h04E4] <= 32'hFED44783;
    mem['h04E5] <= 32'h00278793;
    mem['h04E6] <= 32'h02F71C63;
    mem['h04E7] <= 32'hFEF44703;
    mem['h04E8] <= 32'h00070793;
    mem['h04E9] <= 32'h00279793;
    mem['h04EA] <= 32'h00E787B3;
    mem['h04EB] <= 32'h00379793;
    mem['h04EC] <= 32'h00078713;
    mem['h04ED] <= 32'hFEE44783;
    mem['h04EE] <= 32'h00F707B3;
    mem['h04EF] <= 32'h00279713;
    mem['h04F0] <= 32'h052007B7;
    mem['h04F1] <= 32'h00F707B3;
    mem['h04F2] <= 32'h00200713;
    mem['h04F3] <= 32'h00E7A023;
    mem['h04F4] <= 32'hFEE44703;
    mem['h04F5] <= 32'h01000793;
    mem['h04F6] <= 32'h04F71C63;
    mem['h04F7] <= 32'hFEF44703;
    mem['h04F8] <= 32'hFED44783;
    mem['h04F9] <= 32'h00378793;
    mem['h04FA] <= 32'h00F70A63;
    mem['h04FB] <= 32'hFEF44703;
    mem['h04FC] <= 32'hFED44783;
    mem['h04FD] <= 32'h00478793;
    mem['h04FE] <= 32'h02F71C63;
    mem['h04FF] <= 32'hFEF44703;
    mem['h0500] <= 32'h00070793;
    mem['h0501] <= 32'h00279793;
    mem['h0502] <= 32'h00E787B3;
    mem['h0503] <= 32'h00379793;
    mem['h0504] <= 32'h00078713;
    mem['h0505] <= 32'hFEE44783;
    mem['h0506] <= 32'h00F707B3;
    mem['h0507] <= 32'h00279713;
    mem['h0508] <= 32'h052007B7;
    mem['h0509] <= 32'h00F707B3;
    mem['h050A] <= 32'h00200713;
    mem['h050B] <= 32'h00E7A023;
    mem['h050C] <= 32'hFEE44703;
    mem['h050D] <= 32'h01200793;
    mem['h050E] <= 32'h04F71A63;
    mem['h050F] <= 32'hFEF44703;
    mem['h0510] <= 32'hFED44783;
    mem['h0511] <= 32'h04F76463;
    mem['h0512] <= 32'hFEF44703;
    mem['h0513] <= 32'hFED44783;
    mem['h0514] <= 32'h00478793;
    mem['h0515] <= 32'h02E7CC63;
    mem['h0516] <= 32'hFEF44703;
    mem['h0517] <= 32'h00070793;
    mem['h0518] <= 32'h00279793;
    mem['h0519] <= 32'h00E787B3;
    mem['h051A] <= 32'h00379793;
    mem['h051B] <= 32'h00078713;
    mem['h051C] <= 32'hFEE44783;
    mem['h051D] <= 32'h00F707B3;
    mem['h051E] <= 32'h00279713;
    mem['h051F] <= 32'h052007B7;
    mem['h0520] <= 32'h00F707B3;
    mem['h0521] <= 32'h00200713;
    mem['h0522] <= 32'h00E7A023;
    mem['h0523] <= 32'hFEF44703;
    mem['h0524] <= 32'hFED44783;
    mem['h0525] <= 32'h04F71863;
    mem['h0526] <= 32'hFEE44703;
    mem['h0527] <= 32'h01400793;
    mem['h0528] <= 32'h00F70863;
    mem['h0529] <= 32'hFEE44703;
    mem['h052A] <= 32'h01500793;
    mem['h052B] <= 32'h02F71C63;
    mem['h052C] <= 32'hFEF44703;
    mem['h052D] <= 32'h00070793;
    mem['h052E] <= 32'h00279793;
    mem['h052F] <= 32'h00E787B3;
    mem['h0530] <= 32'h00379793;
    mem['h0531] <= 32'h00078713;
    mem['h0532] <= 32'hFEE44783;
    mem['h0533] <= 32'h00F707B3;
    mem['h0534] <= 32'h00279713;
    mem['h0535] <= 32'h052007B7;
    mem['h0536] <= 32'h00F707B3;
    mem['h0537] <= 32'h00700713;
    mem['h0538] <= 32'h00E7A023;
    mem['h0539] <= 32'hFEE44703;
    mem['h053A] <= 32'h01400793;
    mem['h053B] <= 32'h06F71463;
    mem['h053C] <= 32'hFEF44703;
    mem['h053D] <= 32'hFED44783;
    mem['h053E] <= 32'h00178793;
    mem['h053F] <= 32'h02F70263;
    mem['h0540] <= 32'hFEF44703;
    mem['h0541] <= 32'hFED44783;
    mem['h0542] <= 32'h00278793;
    mem['h0543] <= 32'h00F70A63;
    mem['h0544] <= 32'hFEF44703;
    mem['h0545] <= 32'hFED44783;
    mem['h0546] <= 32'h00478793;
    mem['h0547] <= 32'h02F71C63;
    mem['h0548] <= 32'hFEF44703;
    mem['h0549] <= 32'h00070793;
    mem['h054A] <= 32'h00279793;
    mem['h054B] <= 32'h00E787B3;
    mem['h054C] <= 32'h00379793;
    mem['h054D] <= 32'h00078713;
    mem['h054E] <= 32'hFEE44783;
    mem['h054F] <= 32'h00F707B3;
    mem['h0550] <= 32'h00279713;
    mem['h0551] <= 32'h052007B7;
    mem['h0552] <= 32'h00F707B3;
    mem['h0553] <= 32'h00700713;
    mem['h0554] <= 32'h00E7A023;
    mem['h0555] <= 32'hFEE44703;
    mem['h0556] <= 32'h01500793;
    mem['h0557] <= 32'h04F71C63;
    mem['h0558] <= 32'hFED44783;
    mem['h0559] <= 32'h00178713;
    mem['h055A] <= 32'hFEF44783;
    mem['h055B] <= 32'h04F75463;
    mem['h055C] <= 32'hFEF44703;
    mem['h055D] <= 32'hFED44783;
    mem['h055E] <= 32'h00478793;
    mem['h055F] <= 32'h02E7CC63;
    mem['h0560] <= 32'hFEF44703;
    mem['h0561] <= 32'h00070793;
    mem['h0562] <= 32'h00279793;
    mem['h0563] <= 32'h00E787B3;
    mem['h0564] <= 32'h00379793;
    mem['h0565] <= 32'h00078713;
    mem['h0566] <= 32'hFEE44783;
    mem['h0567] <= 32'h00F707B3;
    mem['h0568] <= 32'h00279713;
    mem['h0569] <= 32'h052007B7;
    mem['h056A] <= 32'h00F707B3;
    mem['h056B] <= 32'h00700713;
    mem['h056C] <= 32'h00E7A023;
    mem['h056D] <= 32'hFEE44703;
    mem['h056E] <= 32'h01700793;
    mem['h056F] <= 32'h00F70863;
    mem['h0570] <= 32'hFEE44703;
    mem['h0571] <= 32'h01900793;
    mem['h0572] <= 32'h04F71A63;
    mem['h0573] <= 32'hFED44703;
    mem['h0574] <= 32'hFEF44783;
    mem['h0575] <= 32'h04F77463;
    mem['h0576] <= 32'hFEF44703;
    mem['h0577] <= 32'hFED44783;
    mem['h0578] <= 32'h00478793;
    mem['h0579] <= 32'h02E7CC63;
    mem['h057A] <= 32'hFEF44703;
    mem['h057B] <= 32'h00070793;
    mem['h057C] <= 32'h00279793;
    mem['h057D] <= 32'h00E787B3;
    mem['h057E] <= 32'h00379793;
    mem['h057F] <= 32'h00078713;
    mem['h0580] <= 32'hFEE44783;
    mem['h0581] <= 32'h00F707B3;
    mem['h0582] <= 32'h00279713;
    mem['h0583] <= 32'h052007B7;
    mem['h0584] <= 32'h00F707B3;
    mem['h0585] <= 32'h00700713;
    mem['h0586] <= 32'h00E7A023;
    mem['h0587] <= 32'hFEE44703;
    mem['h0588] <= 32'h01800793;
    mem['h0589] <= 32'h04F71463;
    mem['h058A] <= 32'hFEF44703;
    mem['h058B] <= 32'hFED44783;
    mem['h058C] <= 32'h00278793;
    mem['h058D] <= 32'h02F71C63;
    mem['h058E] <= 32'hFEF44703;
    mem['h058F] <= 32'h00070793;
    mem['h0590] <= 32'h00279793;
    mem['h0591] <= 32'h00E787B3;
    mem['h0592] <= 32'h00379793;
    mem['h0593] <= 32'h00078713;
    mem['h0594] <= 32'hFEE44783;
    mem['h0595] <= 32'h00F707B3;
    mem['h0596] <= 32'h00279713;
    mem['h0597] <= 32'h052007B7;
    mem['h0598] <= 32'h00F707B3;
    mem['h0599] <= 32'h00700713;
    mem['h059A] <= 32'h00E7A023;
    mem['h059B] <= 32'hFEE44703;
    mem['h059C] <= 32'h01800793;
    mem['h059D] <= 32'h04F71263;
    mem['h059E] <= 32'hFEF44703;
    mem['h059F] <= 32'hFED44783;
    mem['h05A0] <= 32'h02F71C63;
    mem['h05A1] <= 32'hFEF44703;
    mem['h05A2] <= 32'h00070793;
    mem['h05A3] <= 32'h00279793;
    mem['h05A4] <= 32'h00E787B3;
    mem['h05A5] <= 32'h00379793;
    mem['h05A6] <= 32'h00078713;
    mem['h05A7] <= 32'hFEE44783;
    mem['h05A8] <= 32'h00F707B3;
    mem['h05A9] <= 32'h00279713;
    mem['h05AA] <= 32'h052007B7;
    mem['h05AB] <= 32'h00F707B3;
    mem['h05AC] <= 32'h00700713;
    mem['h05AD] <= 32'h00E7A023;
    mem['h05AE] <= 32'hFEE44703;
    mem['h05AF] <= 32'h01B00793;
    mem['h05B0] <= 32'h04F71A63;
    mem['h05B1] <= 32'hFEF44703;
    mem['h05B2] <= 32'hFED44783;
    mem['h05B3] <= 32'h04F76463;
    mem['h05B4] <= 32'hFEF44703;
    mem['h05B5] <= 32'hFED44783;
    mem['h05B6] <= 32'h00478793;
    mem['h05B7] <= 32'h02E7CC63;
    mem['h05B8] <= 32'hFEF44703;
    mem['h05B9] <= 32'h00070793;
    mem['h05BA] <= 32'h00279793;
    mem['h05BB] <= 32'h00E787B3;
    mem['h05BC] <= 32'h00379793;
    mem['h05BD] <= 32'h00078713;
    mem['h05BE] <= 32'hFEE44783;
    mem['h05BF] <= 32'h00F707B3;
    mem['h05C0] <= 32'h00279713;
    mem['h05C1] <= 32'h052007B7;
    mem['h05C2] <= 32'h00F707B3;
    mem['h05C3] <= 32'h00700713;
    mem['h05C4] <= 32'h00E7A023;
    mem['h05C5] <= 32'hFEE44703;
    mem['h05C6] <= 32'h01C00793;
    mem['h05C7] <= 32'h04F71263;
    mem['h05C8] <= 32'hFEF44703;
    mem['h05C9] <= 32'hFED44783;
    mem['h05CA] <= 32'h02F71C63;
    mem['h05CB] <= 32'hFEF44703;
    mem['h05CC] <= 32'h00070793;
    mem['h05CD] <= 32'h00279793;
    mem['h05CE] <= 32'h00E787B3;
    mem['h05CF] <= 32'h00379793;
    mem['h05D0] <= 32'h00078713;
    mem['h05D1] <= 32'hFEE44783;
    mem['h05D2] <= 32'h00F707B3;
    mem['h05D3] <= 32'h00279713;
    mem['h05D4] <= 32'h052007B7;
    mem['h05D5] <= 32'h00F707B3;
    mem['h05D6] <= 32'h00700713;
    mem['h05D7] <= 32'h00E7A023;
    mem['h05D8] <= 32'hFEE44703;
    mem['h05D9] <= 32'h01D00793;
    mem['h05DA] <= 32'h04F71463;
    mem['h05DB] <= 32'hFEF44703;
    mem['h05DC] <= 32'hFED44783;
    mem['h05DD] <= 32'h00178793;
    mem['h05DE] <= 32'h02F71C63;
    mem['h05DF] <= 32'hFEF44703;
    mem['h05E0] <= 32'h00070793;
    mem['h05E1] <= 32'h00279793;
    mem['h05E2] <= 32'h00E787B3;
    mem['h05E3] <= 32'h00379793;
    mem['h05E4] <= 32'h00078713;
    mem['h05E5] <= 32'hFEE44783;
    mem['h05E6] <= 32'h00F707B3;
    mem['h05E7] <= 32'h00279713;
    mem['h05E8] <= 32'h052007B7;
    mem['h05E9] <= 32'h00F707B3;
    mem['h05EA] <= 32'h00700713;
    mem['h05EB] <= 32'h00E7A023;
    mem['h05EC] <= 32'hFEE44703;
    mem['h05ED] <= 32'h01C00793;
    mem['h05EE] <= 32'h04F71463;
    mem['h05EF] <= 32'hFEF44703;
    mem['h05F0] <= 32'hFED44783;
    mem['h05F1] <= 32'h00278793;
    mem['h05F2] <= 32'h02F71C63;
    mem['h05F3] <= 32'hFEF44703;
    mem['h05F4] <= 32'h00070793;
    mem['h05F5] <= 32'h00279793;
    mem['h05F6] <= 32'h00E787B3;
    mem['h05F7] <= 32'h00379793;
    mem['h05F8] <= 32'h00078713;
    mem['h05F9] <= 32'hFEE44783;
    mem['h05FA] <= 32'h00F707B3;
    mem['h05FB] <= 32'h00279713;
    mem['h05FC] <= 32'h052007B7;
    mem['h05FD] <= 32'h00F707B3;
    mem['h05FE] <= 32'h00700713;
    mem['h05FF] <= 32'h00E7A023;
    mem['h0600] <= 32'hFEE44703;
    mem['h0601] <= 32'h01D00793;
    mem['h0602] <= 32'h04F71C63;
    mem['h0603] <= 32'hFEF44703;
    mem['h0604] <= 32'hFED44783;
    mem['h0605] <= 32'h00378793;
    mem['h0606] <= 32'h00F70A63;
    mem['h0607] <= 32'hFEF44703;
    mem['h0608] <= 32'hFED44783;
    mem['h0609] <= 32'h00478793;
    mem['h060A] <= 32'h02F71C63;
    mem['h060B] <= 32'hFEF44703;
    mem['h060C] <= 32'h00070793;
    mem['h060D] <= 32'h00279793;
    mem['h060E] <= 32'h00E787B3;
    mem['h060F] <= 32'h00379793;
    mem['h0610] <= 32'h00078713;
    mem['h0611] <= 32'hFEE44783;
    mem['h0612] <= 32'h00F707B3;
    mem['h0613] <= 32'h00279713;
    mem['h0614] <= 32'h052007B7;
    mem['h0615] <= 32'h00F707B3;
    mem['h0616] <= 32'h00700713;
    mem['h0617] <= 32'h00E7A023;
    mem['h0618] <= 32'hFEE44703;
    mem['h0619] <= 32'h01F00793;
    mem['h061A] <= 32'h00F70863;
    mem['h061B] <= 32'hFEE44703;
    mem['h061C] <= 32'h02100793;
    mem['h061D] <= 32'h04F71A63;
    mem['h061E] <= 32'hFED44703;
    mem['h061F] <= 32'hFEF44783;
    mem['h0620] <= 32'h04F77463;
    mem['h0621] <= 32'hFEF44703;
    mem['h0622] <= 32'hFED44783;
    mem['h0623] <= 32'h00478793;
    mem['h0624] <= 32'h02E7CC63;
    mem['h0625] <= 32'hFEF44703;
    mem['h0626] <= 32'h00070793;
    mem['h0627] <= 32'h00279793;
    mem['h0628] <= 32'h00E787B3;
    mem['h0629] <= 32'h00379793;
    mem['h062A] <= 32'h00078713;
    mem['h062B] <= 32'hFEE44783;
    mem['h062C] <= 32'h00F707B3;
    mem['h062D] <= 32'h00279713;
    mem['h062E] <= 32'h052007B7;
    mem['h062F] <= 32'h00F707B3;
    mem['h0630] <= 32'h00700713;
    mem['h0631] <= 32'h00E7A023;
    mem['h0632] <= 32'hFEE44703;
    mem['h0633] <= 32'h02000793;
    mem['h0634] <= 32'h04F71463;
    mem['h0635] <= 32'hFEF44703;
    mem['h0636] <= 32'hFED44783;
    mem['h0637] <= 32'h00278793;
    mem['h0638] <= 32'h02F71C63;
    mem['h0639] <= 32'hFEF44703;
    mem['h063A] <= 32'h00070793;
    mem['h063B] <= 32'h00279793;
    mem['h063C] <= 32'h00E787B3;
    mem['h063D] <= 32'h00379793;
    mem['h063E] <= 32'h00078713;
    mem['h063F] <= 32'hFEE44783;
    mem['h0640] <= 32'h00F707B3;
    mem['h0641] <= 32'h00279713;
    mem['h0642] <= 32'h052007B7;
    mem['h0643] <= 32'h00F707B3;
    mem['h0644] <= 32'h00700713;
    mem['h0645] <= 32'h00E7A023;
    mem['h0646] <= 32'hFEE44703;
    mem['h0647] <= 32'h02000793;
    mem['h0648] <= 32'h04F71263;
    mem['h0649] <= 32'hFEF44703;
    mem['h064A] <= 32'hFED44783;
    mem['h064B] <= 32'h02F71C63;
    mem['h064C] <= 32'hFEF44703;
    mem['h064D] <= 32'h00070793;
    mem['h064E] <= 32'h00279793;
    mem['h064F] <= 32'h00E787B3;
    mem['h0650] <= 32'h00379793;
    mem['h0651] <= 32'h00078713;
    mem['h0652] <= 32'hFEE44783;
    mem['h0653] <= 32'h00F707B3;
    mem['h0654] <= 32'h00279713;
    mem['h0655] <= 32'h052007B7;
    mem['h0656] <= 32'h00F707B3;
    mem['h0657] <= 32'h00700713;
    mem['h0658] <= 32'h00E7A023;
    mem['h0659] <= 32'hFEE44703;
    mem['h065A] <= 32'h02500793;
    mem['h065B] <= 32'h04F71A63;
    mem['h065C] <= 32'hFEF44703;
    mem['h065D] <= 32'hFED44783;
    mem['h065E] <= 32'h04F76463;
    mem['h065F] <= 32'hFEF44703;
    mem['h0660] <= 32'hFED44783;
    mem['h0661] <= 32'h00478793;
    mem['h0662] <= 32'h02E7CC63;
    mem['h0663] <= 32'hFEF44703;
    mem['h0664] <= 32'h00070793;
    mem['h0665] <= 32'h00279793;
    mem['h0666] <= 32'h00E787B3;
    mem['h0667] <= 32'h00379793;
    mem['h0668] <= 32'h00078713;
    mem['h0669] <= 32'hFEE44783;
    mem['h066A] <= 32'h00F707B3;
    mem['h066B] <= 32'h00279713;
    mem['h066C] <= 32'h052007B7;
    mem['h066D] <= 32'h00F707B3;
    mem['h066E] <= 32'h00700713;
    mem['h066F] <= 32'h00E7A023;
    mem['h0670] <= 32'hFEE44703;
    mem['h0671] <= 32'h02300793;
    mem['h0672] <= 32'h00F70863;
    mem['h0673] <= 32'hFEE44703;
    mem['h0674] <= 32'h02400793;
    mem['h0675] <= 32'h04F71463;
    mem['h0676] <= 32'hFEF44703;
    mem['h0677] <= 32'hFED44783;
    mem['h0678] <= 32'h00478793;
    mem['h0679] <= 32'h02F71C63;
    mem['h067A] <= 32'hFEF44703;
    mem['h067B] <= 32'h00070793;
    mem['h067C] <= 32'h00279793;
    mem['h067D] <= 32'h00E787B3;
    mem['h067E] <= 32'h00379793;
    mem['h067F] <= 32'h00078713;
    mem['h0680] <= 32'hFEE44783;
    mem['h0681] <= 32'h00F707B3;
    mem['h0682] <= 32'h00279713;
    mem['h0683] <= 32'h052007B7;
    mem['h0684] <= 32'h00F707B3;
    mem['h0685] <= 32'h00700713;
    mem['h0686] <= 32'h00E7A023;
    mem['h0687] <= 32'hFEE44703;
    mem['h0688] <= 32'h02300793;
    mem['h0689] <= 32'h04F71463;
    mem['h068A] <= 32'hFEF44703;
    mem['h068B] <= 32'hFED44783;
    mem['h068C] <= 32'h00378793;
    mem['h068D] <= 32'h02F71C63;
    mem['h068E] <= 32'hFEF44703;
    mem['h068F] <= 32'h00070793;
    mem['h0690] <= 32'h00279793;
    mem['h0691] <= 32'h00E787B3;
    mem['h0692] <= 32'h00379793;
    mem['h0693] <= 32'h00078713;
    mem['h0694] <= 32'hFEE44783;
    mem['h0695] <= 32'h00F707B3;
    mem['h0696] <= 32'h00279713;
    mem['h0697] <= 32'h052007B7;
    mem['h0698] <= 32'h00F707B3;
    mem['h0699] <= 32'h00700713;
    mem['h069A] <= 32'h00E7A023;
    mem['h069B] <= 32'hFEE44783;
    mem['h069C] <= 32'h00178793;
    mem['h069D] <= 32'hFEF40723;
    mem['h069E] <= 32'hFEE44703;
    mem['h069F] <= 32'h02700793;
    mem['h06A0] <= 32'hDCE7FC63;
    mem['h06A1] <= 32'hFEF44783;
    mem['h06A2] <= 32'h00178793;
    mem['h06A3] <= 32'hFEF407A3;
    mem['h06A4] <= 32'hFEF44703;
    mem['h06A5] <= 32'h01D00793;
    mem['h06A6] <= 32'hDAE7FC63;
    mem['h06A7] <= 32'h00000013;
    mem['h06A8] <= 32'h00000013;
    mem['h06A9] <= 32'h01C12403;
    mem['h06AA] <= 32'h02010113;
    mem['h06AB] <= 32'h00008067;
    mem['h06AC] <= 32'hFD010113;
    mem['h06AD] <= 32'h02812623;
    mem['h06AE] <= 32'h03010413;
    mem['h06AF] <= 32'hFCA42E23;
    mem['h06B0] <= 32'hFCB42C23;
    mem['h06B1] <= 32'hFCC42A23;
    mem['h06B2] <= 32'hFE042623;
    mem['h06B3] <= 32'h6A80006F;
    mem['h06B4] <= 32'hFE042423;
    mem['h06B5] <= 32'h6880006F;
    mem['h06B6] <= 32'hFDC42783;
    mem['h06B7] <= 32'h00278793;
    mem['h06B8] <= 32'hFE842703;
    mem['h06B9] <= 32'h02F70A63;
    mem['h06BA] <= 32'hFDC42783;
    mem['h06BB] <= 32'h00378793;
    mem['h06BC] <= 32'hFE842703;
    mem['h06BD] <= 32'h02F70263;
    mem['h06BE] <= 32'hFDC42783;
    mem['h06BF] <= 32'h00778793;
    mem['h06C0] <= 32'hFE842703;
    mem['h06C1] <= 32'h00F70A63;
    mem['h06C2] <= 32'hFDC42783;
    mem['h06C3] <= 32'h00878793;
    mem['h06C4] <= 32'hFE842703;
    mem['h06C5] <= 32'h04F71063;
    mem['h06C6] <= 32'hFEC42703;
    mem['h06C7] <= 32'hFD842783;
    mem['h06C8] <= 32'h02F71A63;
    mem['h06C9] <= 32'hFEC42703;
    mem['h06CA] <= 32'h00070793;
    mem['h06CB] <= 32'h00279793;
    mem['h06CC] <= 32'h00E787B3;
    mem['h06CD] <= 32'h00379793;
    mem['h06CE] <= 32'h00078713;
    mem['h06CF] <= 32'hFE842783;
    mem['h06D0] <= 32'h00F707B3;
    mem['h06D1] <= 32'h00279713;
    mem['h06D2] <= 32'h052007B7;
    mem['h06D3] <= 32'h00F707B3;
    mem['h06D4] <= 32'h0007A023;
    mem['h06D5] <= 32'hFDC42783;
    mem['h06D6] <= 32'h00178793;
    mem['h06D7] <= 32'hFE842703;
    mem['h06D8] <= 32'h02F70A63;
    mem['h06D9] <= 32'hFDC42783;
    mem['h06DA] <= 32'h00478793;
    mem['h06DB] <= 32'hFE842703;
    mem['h06DC] <= 32'h02F70263;
    mem['h06DD] <= 32'hFDC42783;
    mem['h06DE] <= 32'h00678793;
    mem['h06DF] <= 32'hFE842703;
    mem['h06E0] <= 32'h00F70A63;
    mem['h06E1] <= 32'hFDC42783;
    mem['h06E2] <= 32'h00978793;
    mem['h06E3] <= 32'hFE842703;
    mem['h06E4] <= 32'h04F71263;
    mem['h06E5] <= 32'hFD842783;
    mem['h06E6] <= 32'h00178793;
    mem['h06E7] <= 32'hFEC42703;
    mem['h06E8] <= 32'h02F71A63;
    mem['h06E9] <= 32'hFEC42703;
    mem['h06EA] <= 32'h00070793;
    mem['h06EB] <= 32'h00279793;
    mem['h06EC] <= 32'h00E787B3;
    mem['h06ED] <= 32'h00379793;
    mem['h06EE] <= 32'h00078713;
    mem['h06EF] <= 32'hFE842783;
    mem['h06F0] <= 32'h00F707B3;
    mem['h06F1] <= 32'h00279713;
    mem['h06F2] <= 32'h052007B7;
    mem['h06F3] <= 32'h00F707B3;
    mem['h06F4] <= 32'h0007A023;
    mem['h06F5] <= 32'hFE842703;
    mem['h06F6] <= 32'hFDC42783;
    mem['h06F7] <= 32'h02F70263;
    mem['h06F8] <= 32'hFDC42783;
    mem['h06F9] <= 32'h00578793;
    mem['h06FA] <= 32'hFE842703;
    mem['h06FB] <= 32'h00F70A63;
    mem['h06FC] <= 32'hFDC42783;
    mem['h06FD] <= 32'h00A78793;
    mem['h06FE] <= 32'hFE842703;
    mem['h06FF] <= 32'h04F71263;
    mem['h0700] <= 32'hFD842783;
    mem['h0701] <= 32'h00278793;
    mem['h0702] <= 32'hFEC42703;
    mem['h0703] <= 32'h02F71A63;
    mem['h0704] <= 32'hFEC42703;
    mem['h0705] <= 32'h00070793;
    mem['h0706] <= 32'h00279793;
    mem['h0707] <= 32'h00E787B3;
    mem['h0708] <= 32'h00379793;
    mem['h0709] <= 32'h00078713;
    mem['h070A] <= 32'hFE842783;
    mem['h070B] <= 32'h00F707B3;
    mem['h070C] <= 32'h00279713;
    mem['h070D] <= 32'h052007B7;
    mem['h070E] <= 32'h00F707B3;
    mem['h070F] <= 32'h0007A023;
    mem['h0710] <= 32'hFE842703;
    mem['h0711] <= 32'hFDC42783;
    mem['h0712] <= 32'h00F70A63;
    mem['h0713] <= 32'hFDC42783;
    mem['h0714] <= 32'h00A78793;
    mem['h0715] <= 32'hFE842703;
    mem['h0716] <= 32'h04F71263;
    mem['h0717] <= 32'hFD842783;
    mem['h0718] <= 32'h00378793;
    mem['h0719] <= 32'hFEC42703;
    mem['h071A] <= 32'h02F71A63;
    mem['h071B] <= 32'hFEC42703;
    mem['h071C] <= 32'h00070793;
    mem['h071D] <= 32'h00279793;
    mem['h071E] <= 32'h00E787B3;
    mem['h071F] <= 32'h00379793;
    mem['h0720] <= 32'h00078713;
    mem['h0721] <= 32'hFE842783;
    mem['h0722] <= 32'h00F707B3;
    mem['h0723] <= 32'h00279713;
    mem['h0724] <= 32'h052007B7;
    mem['h0725] <= 32'h00F707B3;
    mem['h0726] <= 32'h0007A023;
    mem['h0727] <= 32'hFDC42783;
    mem['h0728] <= 32'h00178793;
    mem['h0729] <= 32'hFE842703;
    mem['h072A] <= 32'h00F70A63;
    mem['h072B] <= 32'hFDC42783;
    mem['h072C] <= 32'h00978793;
    mem['h072D] <= 32'hFE842703;
    mem['h072E] <= 32'h04F71263;
    mem['h072F] <= 32'hFD842783;
    mem['h0730] <= 32'h00478793;
    mem['h0731] <= 32'hFEC42703;
    mem['h0732] <= 32'h02F71A63;
    mem['h0733] <= 32'hFEC42703;
    mem['h0734] <= 32'h00070793;
    mem['h0735] <= 32'h00279793;
    mem['h0736] <= 32'h00E787B3;
    mem['h0737] <= 32'h00379793;
    mem['h0738] <= 32'h00078713;
    mem['h0739] <= 32'hFE842783;
    mem['h073A] <= 32'h00F707B3;
    mem['h073B] <= 32'h00279713;
    mem['h073C] <= 32'h052007B7;
    mem['h073D] <= 32'h00F707B3;
    mem['h073E] <= 32'h0007A023;
    mem['h073F] <= 32'hFDC42783;
    mem['h0740] <= 32'h00278793;
    mem['h0741] <= 32'hFE842703;
    mem['h0742] <= 32'h00F70A63;
    mem['h0743] <= 32'hFDC42783;
    mem['h0744] <= 32'h00878793;
    mem['h0745] <= 32'hFE842703;
    mem['h0746] <= 32'h04F71263;
    mem['h0747] <= 32'hFD842783;
    mem['h0748] <= 32'h00578793;
    mem['h0749] <= 32'hFEC42703;
    mem['h074A] <= 32'h02F71A63;
    mem['h074B] <= 32'hFEC42703;
    mem['h074C] <= 32'h00070793;
    mem['h074D] <= 32'h00279793;
    mem['h074E] <= 32'h00E787B3;
    mem['h074F] <= 32'h00379793;
    mem['h0750] <= 32'h00078713;
    mem['h0751] <= 32'hFE842783;
    mem['h0752] <= 32'h00F707B3;
    mem['h0753] <= 32'h00279713;
    mem['h0754] <= 32'h052007B7;
    mem['h0755] <= 32'h00F707B3;
    mem['h0756] <= 32'h0007A023;
    mem['h0757] <= 32'hFDC42783;
    mem['h0758] <= 32'h00378793;
    mem['h0759] <= 32'hFE842703;
    mem['h075A] <= 32'h00F70A63;
    mem['h075B] <= 32'hFDC42783;
    mem['h075C] <= 32'h00778793;
    mem['h075D] <= 32'hFE842703;
    mem['h075E] <= 32'h04F71263;
    mem['h075F] <= 32'hFD842783;
    mem['h0760] <= 32'h00678793;
    mem['h0761] <= 32'hFEC42703;
    mem['h0762] <= 32'h02F71A63;
    mem['h0763] <= 32'hFEC42703;
    mem['h0764] <= 32'h00070793;
    mem['h0765] <= 32'h00279793;
    mem['h0766] <= 32'h00E787B3;
    mem['h0767] <= 32'h00379793;
    mem['h0768] <= 32'h00078713;
    mem['h0769] <= 32'hFE842783;
    mem['h076A] <= 32'h00F707B3;
    mem['h076B] <= 32'h00279713;
    mem['h076C] <= 32'h052007B7;
    mem['h076D] <= 32'h00F707B3;
    mem['h076E] <= 32'h0007A023;
    mem['h076F] <= 32'hFDC42783;
    mem['h0770] <= 32'h00478793;
    mem['h0771] <= 32'hFE842703;
    mem['h0772] <= 32'h00F70A63;
    mem['h0773] <= 32'hFDC42783;
    mem['h0774] <= 32'h00678793;
    mem['h0775] <= 32'hFE842703;
    mem['h0776] <= 32'h04F71263;
    mem['h0777] <= 32'hFD842783;
    mem['h0778] <= 32'h00778793;
    mem['h0779] <= 32'hFEC42703;
    mem['h077A] <= 32'h02F71A63;
    mem['h077B] <= 32'hFEC42703;
    mem['h077C] <= 32'h00070793;
    mem['h077D] <= 32'h00279793;
    mem['h077E] <= 32'h00E787B3;
    mem['h077F] <= 32'h00379793;
    mem['h0780] <= 32'h00078713;
    mem['h0781] <= 32'hFE842783;
    mem['h0782] <= 32'h00F707B3;
    mem['h0783] <= 32'h00279713;
    mem['h0784] <= 32'h052007B7;
    mem['h0785] <= 32'h00F707B3;
    mem['h0786] <= 32'h0007A023;
    mem['h0787] <= 32'hFDC42783;
    mem['h0788] <= 32'h00578793;
    mem['h0789] <= 32'hFE842703;
    mem['h078A] <= 32'h04F71263;
    mem['h078B] <= 32'hFD842783;
    mem['h078C] <= 32'h00878793;
    mem['h078D] <= 32'hFEC42703;
    mem['h078E] <= 32'h02F71A63;
    mem['h078F] <= 32'hFEC42703;
    mem['h0790] <= 32'h00070793;
    mem['h0791] <= 32'h00279793;
    mem['h0792] <= 32'h00E787B3;
    mem['h0793] <= 32'h00379793;
    mem['h0794] <= 32'h00078713;
    mem['h0795] <= 32'hFE842783;
    mem['h0796] <= 32'h00F707B3;
    mem['h0797] <= 32'h00279713;
    mem['h0798] <= 32'h052007B7;
    mem['h0799] <= 32'h00F707B3;
    mem['h079A] <= 32'h0007A023;
    mem['h079B] <= 32'hFDC42783;
    mem['h079C] <= 32'h00278793;
    mem['h079D] <= 32'hFE842703;
    mem['h079E] <= 32'h02F70A63;
    mem['h079F] <= 32'hFDC42783;
    mem['h07A0] <= 32'h00378793;
    mem['h07A1] <= 32'hFE842703;
    mem['h07A2] <= 32'h02F70263;
    mem['h07A3] <= 32'hFDC42783;
    mem['h07A4] <= 32'h00778793;
    mem['h07A5] <= 32'hFE842703;
    mem['h07A6] <= 32'h00F70A63;
    mem['h07A7] <= 32'hFDC42783;
    mem['h07A8] <= 32'h00878793;
    mem['h07A9] <= 32'hFE842703;
    mem['h07AA] <= 32'h04F71463;
    mem['h07AB] <= 32'hFD842783;
    mem['h07AC] <= 32'h00178793;
    mem['h07AD] <= 32'hFEC42703;
    mem['h07AE] <= 32'h02F71C63;
    mem['h07AF] <= 32'hFEC42703;
    mem['h07B0] <= 32'h00070793;
    mem['h07B1] <= 32'h00279793;
    mem['h07B2] <= 32'h00E787B3;
    mem['h07B3] <= 32'h00379793;
    mem['h07B4] <= 32'h00078713;
    mem['h07B5] <= 32'hFE842783;
    mem['h07B6] <= 32'h00F707B3;
    mem['h07B7] <= 32'h00279713;
    mem['h07B8] <= 32'h052007B7;
    mem['h07B9] <= 32'h00F707B3;
    mem['h07BA] <= 32'hFD442703;
    mem['h07BB] <= 32'h00E7A023;
    mem['h07BC] <= 32'hFDC42703;
    mem['h07BD] <= 32'hFE842783;
    mem['h07BE] <= 32'h00F75A63;
    mem['h07BF] <= 32'hFDC42783;
    mem['h07C0] <= 32'h00478793;
    mem['h07C1] <= 32'hFE842703;
    mem['h07C2] <= 32'h02E7D263;
    mem['h07C3] <= 32'hFDC42783;
    mem['h07C4] <= 32'h00578793;
    mem['h07C5] <= 32'hFE842703;
    mem['h07C6] <= 32'h04E7DC63;
    mem['h07C7] <= 32'hFDC42783;
    mem['h07C8] <= 32'h00978793;
    mem['h07C9] <= 32'hFE842703;
    mem['h07CA] <= 32'h04E7C463;
    mem['h07CB] <= 32'hFD842783;
    mem['h07CC] <= 32'h00278793;
    mem['h07CD] <= 32'hFEC42703;
    mem['h07CE] <= 32'h02F71C63;
    mem['h07CF] <= 32'hFEC42703;
    mem['h07D0] <= 32'h00070793;
    mem['h07D1] <= 32'h00279793;
    mem['h07D2] <= 32'h00E787B3;
    mem['h07D3] <= 32'h00379793;
    mem['h07D4] <= 32'h00078713;
    mem['h07D5] <= 32'hFE842783;
    mem['h07D6] <= 32'h00F707B3;
    mem['h07D7] <= 32'h00279713;
    mem['h07D8] <= 32'h052007B7;
    mem['h07D9] <= 32'h00F707B3;
    mem['h07DA] <= 32'hFD442703;
    mem['h07DB] <= 32'h00E7A023;
    mem['h07DC] <= 32'hFDC42703;
    mem['h07DD] <= 32'hFE842783;
    mem['h07DE] <= 32'h04F75C63;
    mem['h07DF] <= 32'hFDC42783;
    mem['h07E0] <= 32'h00978793;
    mem['h07E1] <= 32'hFE842703;
    mem['h07E2] <= 32'h04E7C463;
    mem['h07E3] <= 32'hFD842783;
    mem['h07E4] <= 32'h00378793;
    mem['h07E5] <= 32'hFEC42703;
    mem['h07E6] <= 32'h02F71C63;
    mem['h07E7] <= 32'hFEC42703;
    mem['h07E8] <= 32'h00070793;
    mem['h07E9] <= 32'h00279793;
    mem['h07EA] <= 32'h00E787B3;
    mem['h07EB] <= 32'h00379793;
    mem['h07EC] <= 32'h00078713;
    mem['h07ED] <= 32'hFE842783;
    mem['h07EE] <= 32'h00F707B3;
    mem['h07EF] <= 32'h00279713;
    mem['h07F0] <= 32'h052007B7;
    mem['h07F1] <= 32'h00F707B3;
    mem['h07F2] <= 32'hFD442703;
    mem['h07F3] <= 32'h00E7A023;
    mem['h07F4] <= 32'hFDC42783;
    mem['h07F5] <= 32'h00178793;
    mem['h07F6] <= 32'hFE842703;
    mem['h07F7] <= 32'h04E7DC63;
    mem['h07F8] <= 32'hFDC42783;
    mem['h07F9] <= 32'h00878793;
    mem['h07FA] <= 32'hFE842703;
    mem['h07FB] <= 32'h04E7C463;
    mem['h07FC] <= 32'hFD842783;
    mem['h07FD] <= 32'h00478793;
    mem['h07FE] <= 32'hFEC42703;
    mem['h07FF] <= 32'h02F71C63;
    mem['h0800] <= 32'hFEC42703;
    mem['h0801] <= 32'h00070793;
    mem['h0802] <= 32'h00279793;
    mem['h0803] <= 32'h00E787B3;
    mem['h0804] <= 32'h00379793;
    mem['h0805] <= 32'h00078713;
    mem['h0806] <= 32'hFE842783;
    mem['h0807] <= 32'h00F707B3;
    mem['h0808] <= 32'h00279713;
    mem['h0809] <= 32'h052007B7;
    mem['h080A] <= 32'h00F707B3;
    mem['h080B] <= 32'hFD442703;
    mem['h080C] <= 32'h00E7A023;
    mem['h080D] <= 32'hFDC42783;
    mem['h080E] <= 32'h00278793;
    mem['h080F] <= 32'hFE842703;
    mem['h0810] <= 32'h04E7DC63;
    mem['h0811] <= 32'hFDC42783;
    mem['h0812] <= 32'h00778793;
    mem['h0813] <= 32'hFE842703;
    mem['h0814] <= 32'h04E7C463;
    mem['h0815] <= 32'hFD842783;
    mem['h0816] <= 32'h00578793;
    mem['h0817] <= 32'hFEC42703;
    mem['h0818] <= 32'h02F71C63;
    mem['h0819] <= 32'hFEC42703;
    mem['h081A] <= 32'h00070793;
    mem['h081B] <= 32'h00279793;
    mem['h081C] <= 32'h00E787B3;
    mem['h081D] <= 32'h00379793;
    mem['h081E] <= 32'h00078713;
    mem['h081F] <= 32'hFE842783;
    mem['h0820] <= 32'h00F707B3;
    mem['h0821] <= 32'h00279713;
    mem['h0822] <= 32'h052007B7;
    mem['h0823] <= 32'h00F707B3;
    mem['h0824] <= 32'hFD442703;
    mem['h0825] <= 32'h00E7A023;
    mem['h0826] <= 32'hFDC42783;
    mem['h0827] <= 32'h00378793;
    mem['h0828] <= 32'hFE842703;
    mem['h0829] <= 32'h04E7DC63;
    mem['h082A] <= 32'hFDC42783;
    mem['h082B] <= 32'h00678793;
    mem['h082C] <= 32'hFE842703;
    mem['h082D] <= 32'h04E7C463;
    mem['h082E] <= 32'hFD842783;
    mem['h082F] <= 32'h00678793;
    mem['h0830] <= 32'hFEC42703;
    mem['h0831] <= 32'h02F71C63;
    mem['h0832] <= 32'hFEC42703;
    mem['h0833] <= 32'h00070793;
    mem['h0834] <= 32'h00279793;
    mem['h0835] <= 32'h00E787B3;
    mem['h0836] <= 32'h00379793;
    mem['h0837] <= 32'h00078713;
    mem['h0838] <= 32'hFE842783;
    mem['h0839] <= 32'h00F707B3;
    mem['h083A] <= 32'h00279713;
    mem['h083B] <= 32'h052007B7;
    mem['h083C] <= 32'h00F707B3;
    mem['h083D] <= 32'hFD442703;
    mem['h083E] <= 32'h00E7A023;
    mem['h083F] <= 32'hFDC42783;
    mem['h0840] <= 32'h00578793;
    mem['h0841] <= 32'hFE842703;
    mem['h0842] <= 32'h04F71463;
    mem['h0843] <= 32'hFD842783;
    mem['h0844] <= 32'h00778793;
    mem['h0845] <= 32'hFEC42703;
    mem['h0846] <= 32'h02F71C63;
    mem['h0847] <= 32'hFEC42703;
    mem['h0848] <= 32'h00070793;
    mem['h0849] <= 32'h00279793;
    mem['h084A] <= 32'h00E787B3;
    mem['h084B] <= 32'h00379793;
    mem['h084C] <= 32'h00078713;
    mem['h084D] <= 32'hFE842783;
    mem['h084E] <= 32'h00F707B3;
    mem['h084F] <= 32'h00279713;
    mem['h0850] <= 32'h052007B7;
    mem['h0851] <= 32'h00F707B3;
    mem['h0852] <= 32'hFD442703;
    mem['h0853] <= 32'h00E7A023;
    mem['h0854] <= 32'hFE842783;
    mem['h0855] <= 32'h00178793;
    mem['h0856] <= 32'hFEF42423;
    mem['h0857] <= 32'hFE842703;
    mem['h0858] <= 32'h02700793;
    mem['h0859] <= 32'h96E7DAE3;
    mem['h085A] <= 32'hFEC42783;
    mem['h085B] <= 32'h00178793;
    mem['h085C] <= 32'hFEF42623;
    mem['h085D] <= 32'hFEC42703;
    mem['h085E] <= 32'h01D00793;
    mem['h085F] <= 32'h94E7DAE3;
    mem['h0860] <= 32'h00000013;
    mem['h0861] <= 32'h00000013;
    mem['h0862] <= 32'h02C12403;
    mem['h0863] <= 32'h03010113;
    mem['h0864] <= 32'h00008067;
    mem['h0865] <= 32'hFD010113;
    mem['h0866] <= 32'h02812623;
    mem['h0867] <= 32'h03010413;
    mem['h0868] <= 32'hFCA42E23;
    mem['h0869] <= 32'hFE0407A3;
    mem['h086A] <= 32'h0640006F;
    mem['h086B] <= 32'hFE040723;
    mem['h086C] <= 32'h0440006F;
    mem['h086D] <= 32'hFEF44703;
    mem['h086E] <= 32'h00070793;
    mem['h086F] <= 32'h00279793;
    mem['h0870] <= 32'h00E787B3;
    mem['h0871] <= 32'h00379793;
    mem['h0872] <= 32'h00078713;
    mem['h0873] <= 32'hFEE44783;
    mem['h0874] <= 32'h00F707B3;
    mem['h0875] <= 32'h00279713;
    mem['h0876] <= 32'h052007B7;
    mem['h0877] <= 32'h00F707B3;
    mem['h0878] <= 32'hFDC42703;
    mem['h0879] <= 32'h00E7A023;
    mem['h087A] <= 32'hFEE44783;
    mem['h087B] <= 32'h00178793;
    mem['h087C] <= 32'hFEF40723;
    mem['h087D] <= 32'hFEE44703;
    mem['h087E] <= 32'h02700793;
    mem['h087F] <= 32'hFAE7FCE3;
    mem['h0880] <= 32'hFEF44783;
    mem['h0881] <= 32'h00178793;
    mem['h0882] <= 32'hFEF407A3;
    mem['h0883] <= 32'hFEF44703;
    mem['h0884] <= 32'h01D00793;
    mem['h0885] <= 32'hF8E7FCE3;
    mem['h0886] <= 32'h00000013;
    mem['h0887] <= 32'h00000013;
    mem['h0888] <= 32'h02C12403;
    mem['h0889] <= 32'h03010113;
    mem['h088A] <= 32'h00008067;
    mem['h088B] <= 32'hFD010113;
    mem['h088C] <= 32'h02112623;
    mem['h088D] <= 32'h02812423;
    mem['h088E] <= 32'h03010413;
    mem['h088F] <= 32'hFCA42E23;
    mem['h0890] <= 32'h00100793;
    mem['h0891] <= 32'hFEF406A3;
    mem['h0892] <= 32'hFE0407A3;
    mem['h0893] <= 32'h7980006F;
    mem['h0894] <= 32'hFE040723;
    mem['h0895] <= 32'h7780006F;
    mem['h0896] <= 32'hFEF44703;
    mem['h0897] <= 32'h00070793;
    mem['h0898] <= 32'h00279793;
    mem['h0899] <= 32'h00E787B3;
    mem['h089A] <= 32'h00379793;
    mem['h089B] <= 32'h00078713;
    mem['h089C] <= 32'hFEE44783;
    mem['h089D] <= 32'h00F707B3;
    mem['h089E] <= 32'h00279713;
    mem['h089F] <= 32'h052007B7;
    mem['h08A0] <= 32'h00F707B3;
    mem['h08A1] <= 32'h00900713;
    mem['h08A2] <= 32'h00E7A023;
    mem['h08A3] <= 32'hFEE44703;
    mem['h08A4] <= 32'h00500793;
    mem['h08A5] <= 32'h02F71263;
    mem['h08A6] <= 32'hFED44783;
    mem['h08A7] <= 32'h00178713;
    mem['h08A8] <= 32'hFEF44783;
    mem['h08A9] <= 32'h00F75A63;
    mem['h08AA] <= 32'hFEF44703;
    mem['h08AB] <= 32'hFED44783;
    mem['h08AC] <= 32'h00578793;
    mem['h08AD] <= 32'h0AE7DC63;
    mem['h08AE] <= 32'hFEE44703;
    mem['h08AF] <= 32'h00600793;
    mem['h08B0] <= 32'h02F71263;
    mem['h08B1] <= 32'hFEF44703;
    mem['h08B2] <= 32'hFED44783;
    mem['h08B3] <= 32'h00178793;
    mem['h08B4] <= 32'h08F70E63;
    mem['h08B5] <= 32'hFEF44703;
    mem['h08B6] <= 32'hFED44783;
    mem['h08B7] <= 32'h00678793;
    mem['h08B8] <= 32'h08F70663;
    mem['h08B9] <= 32'hFEE44703;
    mem['h08BA] <= 32'h00600793;
    mem['h08BB] <= 32'h02E7F663;
    mem['h08BC] <= 32'hFEE44703;
    mem['h08BD] <= 32'h00B00793;
    mem['h08BE] <= 32'h02E7E063;
    mem['h08BF] <= 32'hFEF44703;
    mem['h08C0] <= 32'hFED44783;
    mem['h08C1] <= 32'h06F70463;
    mem['h08C2] <= 32'hFEF44703;
    mem['h08C3] <= 32'hFED44783;
    mem['h08C4] <= 32'h00778793;
    mem['h08C5] <= 32'h04F70C63;
    mem['h08C6] <= 32'hFEE44703;
    mem['h08C7] <= 32'h00B00793;
    mem['h08C8] <= 32'h02F71263;
    mem['h08C9] <= 32'hFED44783;
    mem['h08CA] <= 32'h00378713;
    mem['h08CB] <= 32'hFEF44783;
    mem['h08CC] <= 32'h00F75A63;
    mem['h08CD] <= 32'hFEF44703;
    mem['h08CE] <= 32'hFED44783;
    mem['h08CF] <= 32'h00778793;
    mem['h08D0] <= 32'h02E7D663;
    mem['h08D1] <= 32'hFEE44703;
    mem['h08D2] <= 32'h00700793;
    mem['h08D3] <= 32'h04E7FA63;
    mem['h08D4] <= 32'hFEE44703;
    mem['h08D5] <= 32'h00B00793;
    mem['h08D6] <= 32'h04E7E463;
    mem['h08D7] <= 32'hFEF44703;
    mem['h08D8] <= 32'hFED44783;
    mem['h08D9] <= 32'h00478793;
    mem['h08DA] <= 32'h02F71C63;
    mem['h08DB] <= 32'hFEF44703;
    mem['h08DC] <= 32'h00070793;
    mem['h08DD] <= 32'h00279793;
    mem['h08DE] <= 32'h00E787B3;
    mem['h08DF] <= 32'h00379793;
    mem['h08E0] <= 32'h00078713;
    mem['h08E1] <= 32'hFEE44783;
    mem['h08E2] <= 32'h00F707B3;
    mem['h08E3] <= 32'h00279713;
    mem['h08E4] <= 32'h052007B7;
    mem['h08E5] <= 32'h00F707B3;
    mem['h08E6] <= 32'h00300713;
    mem['h08E7] <= 32'h00E7A023;
    mem['h08E8] <= 32'hFEE44703;
    mem['h08E9] <= 32'h01000793;
    mem['h08EA] <= 32'h00F71863;
    mem['h08EB] <= 32'hFEF44703;
    mem['h08EC] <= 32'hFED44783;
    mem['h08ED] <= 32'h0CF70263;
    mem['h08EE] <= 32'hFEE44703;
    mem['h08EF] <= 32'h00F00793;
    mem['h08F0] <= 32'h00F70863;
    mem['h08F1] <= 32'hFEE44703;
    mem['h08F2] <= 32'h01100793;
    mem['h08F3] <= 32'h00F71A63;
    mem['h08F4] <= 32'hFEF44703;
    mem['h08F5] <= 32'hFED44783;
    mem['h08F6] <= 32'h00178793;
    mem['h08F7] <= 32'h08F70E63;
    mem['h08F8] <= 32'hFEE44703;
    mem['h08F9] <= 32'h00E00793;
    mem['h08FA] <= 32'h00F70863;
    mem['h08FB] <= 32'hFEE44703;
    mem['h08FC] <= 32'h01200793;
    mem['h08FD] <= 32'h02F71263;
    mem['h08FE] <= 32'hFED44783;
    mem['h08FF] <= 32'h00178713;
    mem['h0900] <= 32'hFEF44783;
    mem['h0901] <= 32'h00F75A63;
    mem['h0902] <= 32'hFEF44703;
    mem['h0903] <= 32'hFED44783;
    mem['h0904] <= 32'h00378793;
    mem['h0905] <= 32'h06E7D263;
    mem['h0906] <= 32'hFEE44703;
    mem['h0907] <= 32'h00C00793;
    mem['h0908] <= 32'h02E7F063;
    mem['h0909] <= 32'hFEE44703;
    mem['h090A] <= 32'h01300793;
    mem['h090B] <= 32'h00E7EA63;
    mem['h090C] <= 32'hFEF44703;
    mem['h090D] <= 32'hFED44783;
    mem['h090E] <= 32'h00478793;
    mem['h090F] <= 32'h02F70E63;
    mem['h0910] <= 32'hFEE44703;
    mem['h0911] <= 32'h00D00793;
    mem['h0912] <= 32'h00F70863;
    mem['h0913] <= 32'hFEE44703;
    mem['h0914] <= 32'h01300793;
    mem['h0915] <= 32'h04F71C63;
    mem['h0916] <= 32'hFED44783;
    mem['h0917] <= 32'h00478713;
    mem['h0918] <= 32'hFEF44783;
    mem['h0919] <= 32'h04F75463;
    mem['h091A] <= 32'hFEF44703;
    mem['h091B] <= 32'hFED44783;
    mem['h091C] <= 32'h00778793;
    mem['h091D] <= 32'h02E7CC63;
    mem['h091E] <= 32'hFEF44703;
    mem['h091F] <= 32'h00070793;
    mem['h0920] <= 32'h00279793;
    mem['h0921] <= 32'h00E787B3;
    mem['h0922] <= 32'h00379793;
    mem['h0923] <= 32'h00078713;
    mem['h0924] <= 32'hFEE44783;
    mem['h0925] <= 32'h00F707B3;
    mem['h0926] <= 32'h00279713;
    mem['h0927] <= 32'h052007B7;
    mem['h0928] <= 32'h00F707B3;
    mem['h0929] <= 32'h00100713;
    mem['h092A] <= 32'h00E7A023;
    mem['h092B] <= 32'hFEE44703;
    mem['h092C] <= 32'h01500793;
    mem['h092D] <= 32'h00F70863;
    mem['h092E] <= 32'hFEE44703;
    mem['h092F] <= 32'h01C00793;
    mem['h0930] <= 32'h02F71063;
    mem['h0931] <= 32'hFEF44703;
    mem['h0932] <= 32'hFED44783;
    mem['h0933] <= 32'h00F76A63;
    mem['h0934] <= 32'hFEF44703;
    mem['h0935] <= 32'hFED44783;
    mem['h0936] <= 32'h00778793;
    mem['h0937] <= 32'h08E7D263;
    mem['h0938] <= 32'hFEE44703;
    mem['h0939] <= 32'h01600793;
    mem['h093A] <= 32'h00F70863;
    mem['h093B] <= 32'hFEE44703;
    mem['h093C] <= 32'h01B00793;
    mem['h093D] <= 32'h00F71863;
    mem['h093E] <= 32'hFEF44703;
    mem['h093F] <= 32'hFED44783;
    mem['h0940] <= 32'h06F70063;
    mem['h0941] <= 32'hFEE44703;
    mem['h0942] <= 32'h01700793;
    mem['h0943] <= 32'h00F70863;
    mem['h0944] <= 32'hFEE44703;
    mem['h0945] <= 32'h01A00793;
    mem['h0946] <= 32'h02F71063;
    mem['h0947] <= 32'hFED44703;
    mem['h0948] <= 32'hFEF44783;
    mem['h0949] <= 32'h00F77A63;
    mem['h094A] <= 32'hFEF44703;
    mem['h094B] <= 32'hFED44783;
    mem['h094C] <= 32'h00278793;
    mem['h094D] <= 32'h02E7D663;
    mem['h094E] <= 32'hFEE44703;
    mem['h094F] <= 32'h01800793;
    mem['h0950] <= 32'h00F70863;
    mem['h0951] <= 32'hFEE44703;
    mem['h0952] <= 32'h01900793;
    mem['h0953] <= 32'h04F71463;
    mem['h0954] <= 32'hFEF44703;
    mem['h0955] <= 32'hFED44783;
    mem['h0956] <= 32'h00378793;
    mem['h0957] <= 32'h02F71C63;
    mem['h0958] <= 32'hFEF44703;
    mem['h0959] <= 32'h00070793;
    mem['h095A] <= 32'h00279793;
    mem['h095B] <= 32'h00E787B3;
    mem['h095C] <= 32'h00379793;
    mem['h095D] <= 32'h00078713;
    mem['h095E] <= 32'hFEE44783;
    mem['h095F] <= 32'h00F707B3;
    mem['h0960] <= 32'h00279713;
    mem['h0961] <= 32'h052007B7;
    mem['h0962] <= 32'h00F707B3;
    mem['h0963] <= 32'h00200713;
    mem['h0964] <= 32'h00E7A023;
    mem['h0965] <= 32'hFEE44703;
    mem['h0966] <= 32'h01D00793;
    mem['h0967] <= 32'h02E7F663;
    mem['h0968] <= 32'hFEE44703;
    mem['h0969] <= 32'h02200793;
    mem['h096A] <= 32'h02E7E063;
    mem['h096B] <= 32'hFEF44703;
    mem['h096C] <= 32'hFED44783;
    mem['h096D] <= 32'h06F70263;
    mem['h096E] <= 32'hFEF44703;
    mem['h096F] <= 32'hFED44783;
    mem['h0970] <= 32'h00778793;
    mem['h0971] <= 32'h04F70A63;
    mem['h0972] <= 32'hFEE44703;
    mem['h0973] <= 32'h01E00793;
    mem['h0974] <= 32'h02F71063;
    mem['h0975] <= 32'hFED44703;
    mem['h0976] <= 32'hFEF44783;
    mem['h0977] <= 32'h00F77A63;
    mem['h0978] <= 32'hFEF44703;
    mem['h0979] <= 32'hFED44783;
    mem['h097A] <= 32'h00678793;
    mem['h097B] <= 32'h02E7D663;
    mem['h097C] <= 32'hFEE44703;
    mem['h097D] <= 32'h01E00793;
    mem['h097E] <= 32'h04E7FA63;
    mem['h097F] <= 32'hFEE44703;
    mem['h0980] <= 32'h02100793;
    mem['h0981] <= 32'h04E7E463;
    mem['h0982] <= 32'hFEF44703;
    mem['h0983] <= 32'hFED44783;
    mem['h0984] <= 32'h00478793;
    mem['h0985] <= 32'h02F71C63;
    mem['h0986] <= 32'hFEF44703;
    mem['h0987] <= 32'h00070793;
    mem['h0988] <= 32'h00279793;
    mem['h0989] <= 32'h00E787B3;
    mem['h098A] <= 32'h00379793;
    mem['h098B] <= 32'h00078713;
    mem['h098C] <= 32'hFEE44783;
    mem['h098D] <= 32'h00F707B3;
    mem['h098E] <= 32'h00279713;
    mem['h098F] <= 32'h052007B7;
    mem['h0990] <= 32'h00F707B3;
    mem['h0991] <= 32'h00400713;
    mem['h0992] <= 32'h00E7A023;
    mem['h0993] <= 32'hFEE44703;
    mem['h0994] <= 32'h00700793;
    mem['h0995] <= 32'h00F70863;
    mem['h0996] <= 32'hFEE44703;
    mem['h0997] <= 32'h00C00793;
    mem['h0998] <= 32'h02F71263;
    mem['h0999] <= 32'hFED44783;
    mem['h099A] <= 32'h00A78713;
    mem['h099B] <= 32'hFEF44783;
    mem['h099C] <= 32'h00F75A63;
    mem['h099D] <= 32'hFEF44703;
    mem['h099E] <= 32'hFED44783;
    mem['h099F] <= 32'h01078793;
    mem['h09A0] <= 32'h02E7DE63;
    mem['h09A1] <= 32'hFEF44703;
    mem['h09A2] <= 32'hFED44783;
    mem['h09A3] <= 32'h00A78793;
    mem['h09A4] <= 32'h00F70A63;
    mem['h09A5] <= 32'hFEF44703;
    mem['h09A6] <= 32'hFED44783;
    mem['h09A7] <= 32'h01178793;
    mem['h09A8] <= 32'h04F71863;
    mem['h09A9] <= 32'hFEE44703;
    mem['h09AA] <= 32'h00700793;
    mem['h09AB] <= 32'h04E7F263;
    mem['h09AC] <= 32'hFEE44703;
    mem['h09AD] <= 32'h00B00793;
    mem['h09AE] <= 32'h02E7EC63;
    mem['h09AF] <= 32'hFEF44703;
    mem['h09B0] <= 32'h00070793;
    mem['h09B1] <= 32'h00279793;
    mem['h09B2] <= 32'h00E787B3;
    mem['h09B3] <= 32'h00379793;
    mem['h09B4] <= 32'h00078713;
    mem['h09B5] <= 32'hFEE44783;
    mem['h09B6] <= 32'h00F707B3;
    mem['h09B7] <= 32'h00279713;
    mem['h09B8] <= 32'h052007B7;
    mem['h09B9] <= 32'h00F707B3;
    mem['h09BA] <= 32'h00300713;
    mem['h09BB] <= 32'h00E7A023;
    mem['h09BC] <= 32'hFEE44703;
    mem['h09BD] <= 32'h00E00793;
    mem['h09BE] <= 32'h00F70863;
    mem['h09BF] <= 32'hFEE44703;
    mem['h09C0] <= 32'h01400793;
    mem['h09C1] <= 32'h02F71263;
    mem['h09C2] <= 32'hFED44783;
    mem['h09C3] <= 32'h00978713;
    mem['h09C4] <= 32'hFEF44783;
    mem['h09C5] <= 32'h00F75A63;
    mem['h09C6] <= 32'hFEF44703;
    mem['h09C7] <= 32'hFED44783;
    mem['h09C8] <= 32'h00C78793;
    mem['h09C9] <= 32'h08E7D863;
    mem['h09CA] <= 32'hFEE44703;
    mem['h09CB] <= 32'h00F00793;
    mem['h09CC] <= 32'h00F70863;
    mem['h09CD] <= 32'hFEE44703;
    mem['h09CE] <= 32'h01300793;
    mem['h09CF] <= 32'h02F71263;
    mem['h09D0] <= 32'hFED44783;
    mem['h09D1] <= 32'h00C78713;
    mem['h09D2] <= 32'hFEF44783;
    mem['h09D3] <= 32'h00F75A63;
    mem['h09D4] <= 32'hFEF44703;
    mem['h09D5] <= 32'hFED44783;
    mem['h09D6] <= 32'h00E78793;
    mem['h09D7] <= 32'h04E7DC63;
    mem['h09D8] <= 32'hFEE44703;
    mem['h09D9] <= 32'h01000793;
    mem['h09DA] <= 32'h00F70863;
    mem['h09DB] <= 32'hFEE44703;
    mem['h09DC] <= 32'h01200793;
    mem['h09DD] <= 32'h00F71A63;
    mem['h09DE] <= 32'hFEF44703;
    mem['h09DF] <= 32'hFED44783;
    mem['h09E0] <= 32'h00F78793;
    mem['h09E1] <= 32'h02F70863;
    mem['h09E2] <= 32'hFEE44703;
    mem['h09E3] <= 32'h01100793;
    mem['h09E4] <= 32'h04F71C63;
    mem['h09E5] <= 32'hFED44783;
    mem['h09E6] <= 32'h00F78713;
    mem['h09E7] <= 32'hFEF44783;
    mem['h09E8] <= 32'h04F75463;
    mem['h09E9] <= 32'hFEF44703;
    mem['h09EA] <= 32'hFED44783;
    mem['h09EB] <= 32'h01178793;
    mem['h09EC] <= 32'h02E7CC63;
    mem['h09ED] <= 32'hFEF44703;
    mem['h09EE] <= 32'h00070793;
    mem['h09EF] <= 32'h00279793;
    mem['h09F0] <= 32'h00E787B3;
    mem['h09F1] <= 32'h00379793;
    mem['h09F2] <= 32'h00078713;
    mem['h09F3] <= 32'hFEE44783;
    mem['h09F4] <= 32'h00F707B3;
    mem['h09F5] <= 32'h00279713;
    mem['h09F6] <= 32'h052007B7;
    mem['h09F7] <= 32'h00F707B3;
    mem['h09F8] <= 32'h00100713;
    mem['h09F9] <= 32'h00E7A023;
    mem['h09FA] <= 32'hFEE44703;
    mem['h09FB] <= 32'h01500793;
    mem['h09FC] <= 32'h02E7F863;
    mem['h09FD] <= 32'hFEE44703;
    mem['h09FE] <= 32'h01A00793;
    mem['h09FF] <= 32'h02E7E263;
    mem['h0A00] <= 32'hFEF44703;
    mem['h0A01] <= 32'hFED44783;
    mem['h0A02] <= 32'h00A78793;
    mem['h0A03] <= 32'h06F70463;
    mem['h0A04] <= 32'hFEF44703;
    mem['h0A05] <= 32'hFED44783;
    mem['h0A06] <= 32'h01178793;
    mem['h0A07] <= 32'h04F70C63;
    mem['h0A08] <= 32'hFEE44703;
    mem['h0A09] <= 32'h01600793;
    mem['h0A0A] <= 32'h02F71263;
    mem['h0A0B] <= 32'hFED44783;
    mem['h0A0C] <= 32'h00A78713;
    mem['h0A0D] <= 32'hFEF44783;
    mem['h0A0E] <= 32'h00F75A63;
    mem['h0A0F] <= 32'hFEF44703;
    mem['h0A10] <= 32'hFED44783;
    mem['h0A11] <= 32'h01078793;
    mem['h0A12] <= 32'h02E7D663;
    mem['h0A13] <= 32'hFEE44703;
    mem['h0A14] <= 32'h01600793;
    mem['h0A15] <= 32'h04E7FA63;
    mem['h0A16] <= 32'hFEE44703;
    mem['h0A17] <= 32'h01900793;
    mem['h0A18] <= 32'h04E7E463;
    mem['h0A19] <= 32'hFEF44703;
    mem['h0A1A] <= 32'hFED44783;
    mem['h0A1B] <= 32'h00E78793;
    mem['h0A1C] <= 32'h02F71C63;
    mem['h0A1D] <= 32'hFEF44703;
    mem['h0A1E] <= 32'h00070793;
    mem['h0A1F] <= 32'h00279793;
    mem['h0A20] <= 32'h00E787B3;
    mem['h0A21] <= 32'h00379793;
    mem['h0A22] <= 32'h00078713;
    mem['h0A23] <= 32'hFEE44783;
    mem['h0A24] <= 32'h00F707B3;
    mem['h0A25] <= 32'h00279713;
    mem['h0A26] <= 32'h052007B7;
    mem['h0A27] <= 32'h00F707B3;
    mem['h0A28] <= 32'h00200713;
    mem['h0A29] <= 32'h00E7A023;
    mem['h0A2A] <= 32'hFEE44703;
    mem['h0A2B] <= 32'h01C00793;
    mem['h0A2C] <= 32'h02F71263;
    mem['h0A2D] <= 32'hFED44783;
    mem['h0A2E] <= 32'h00978713;
    mem['h0A2F] <= 32'hFEF44783;
    mem['h0A30] <= 32'h00F75A63;
    mem['h0A31] <= 32'hFEF44703;
    mem['h0A32] <= 32'hFED44783;
    mem['h0A33] <= 32'h01178793;
    mem['h0A34] <= 32'h0AE7DE63;
    mem['h0A35] <= 32'hFEE44703;
    mem['h0A36] <= 32'h01C00793;
    mem['h0A37] <= 32'h02E7F863;
    mem['h0A38] <= 32'hFEE44703;
    mem['h0A39] <= 32'h01F00793;
    mem['h0A3A] <= 32'h02E7E263;
    mem['h0A3B] <= 32'hFEF44703;
    mem['h0A3C] <= 32'hFED44783;
    mem['h0A3D] <= 32'h00E78793;
    mem['h0A3E] <= 32'h08F70A63;
    mem['h0A3F] <= 32'hFEF44703;
    mem['h0A40] <= 32'hFED44783;
    mem['h0A41] <= 32'h00A78793;
    mem['h0A42] <= 32'h08F70263;
    mem['h0A43] <= 32'hFEE44703;
    mem['h0A44] <= 32'h02000793;
    mem['h0A45] <= 32'h02F71263;
    mem['h0A46] <= 32'hFED44783;
    mem['h0A47] <= 32'h00A78713;
    mem['h0A48] <= 32'hFEF44783;
    mem['h0A49] <= 32'h00F75A63;
    mem['h0A4A] <= 32'hFEF44703;
    mem['h0A4B] <= 32'hFED44783;
    mem['h0A4C] <= 32'h00D78793;
    mem['h0A4D] <= 32'h04E7DC63;
    mem['h0A4E] <= 32'hFEE44703;
    mem['h0A4F] <= 32'h01E00793;
    mem['h0A50] <= 32'h00F71A63;
    mem['h0A51] <= 32'hFEF44703;
    mem['h0A52] <= 32'hFED44783;
    mem['h0A53] <= 32'h00F78793;
    mem['h0A54] <= 32'h02F70E63;
    mem['h0A55] <= 32'hFEE44703;
    mem['h0A56] <= 32'h01F00793;
    mem['h0A57] <= 32'h00F71A63;
    mem['h0A58] <= 32'hFEF44703;
    mem['h0A59] <= 32'hFED44783;
    mem['h0A5A] <= 32'h01078793;
    mem['h0A5B] <= 32'h02F70063;
    mem['h0A5C] <= 32'hFEE44703;
    mem['h0A5D] <= 32'h02000793;
    mem['h0A5E] <= 32'h04F71463;
    mem['h0A5F] <= 32'hFEF44703;
    mem['h0A60] <= 32'hFED44783;
    mem['h0A61] <= 32'h01178793;
    mem['h0A62] <= 32'h02F71C63;
    mem['h0A63] <= 32'hFEF44703;
    mem['h0A64] <= 32'h00070793;
    mem['h0A65] <= 32'h00279793;
    mem['h0A66] <= 32'h00E787B3;
    mem['h0A67] <= 32'h00379793;
    mem['h0A68] <= 32'h00078713;
    mem['h0A69] <= 32'hFEE44783;
    mem['h0A6A] <= 32'h00F707B3;
    mem['h0A6B] <= 32'h00279713;
    mem['h0A6C] <= 32'h052007B7;
    mem['h0A6D] <= 32'h00F707B3;
    mem['h0A6E] <= 32'h00400713;
    mem['h0A6F] <= 32'h00E7A023;
    mem['h0A70] <= 32'hFEE44783;
    mem['h0A71] <= 32'h00178793;
    mem['h0A72] <= 32'hFEF40723;
    mem['h0A73] <= 32'hFEE44703;
    mem['h0A74] <= 32'h02700793;
    mem['h0A75] <= 32'h88E7F2E3;
    mem['h0A76] <= 32'hFEF44783;
    mem['h0A77] <= 32'h00178793;
    mem['h0A78] <= 32'hFEF407A3;
    mem['h0A79] <= 32'hFEF44703;
    mem['h0A7A] <= 32'h01D00793;
    mem['h0A7B] <= 32'h86E7F2E3;
    mem['h0A7C] <= 32'hFDC42703;
    mem['h0A7D] <= 32'h00300793;
    mem['h0A7E] <= 32'h02F71A63;
    mem['h0A7F] <= 32'h00300613;
    mem['h0A80] <= 32'h01500593;
    mem['h0A81] <= 32'h00500513;
    mem['h0A82] <= 32'h8A8FF0EF;
    mem['h0A83] <= 32'h00300613;
    mem['h0A84] <= 32'h01500593;
    mem['h0A85] <= 32'h00F00513;
    mem['h0A86] <= 32'h898FF0EF;
    mem['h0A87] <= 32'h00300613;
    mem['h0A88] <= 32'h01500593;
    mem['h0A89] <= 32'h01900513;
    mem['h0A8A] <= 32'h888FF0EF;
    mem['h0A8B] <= 32'hFDC42703;
    mem['h0A8C] <= 32'h00200793;
    mem['h0A8D] <= 32'h02F71A63;
    mem['h0A8E] <= 32'h00300613;
    mem['h0A8F] <= 32'h01500593;
    mem['h0A90] <= 32'h00500513;
    mem['h0A91] <= 32'h86CFF0EF;
    mem['h0A92] <= 32'h00300613;
    mem['h0A93] <= 32'h01500593;
    mem['h0A94] <= 32'h00F00513;
    mem['h0A95] <= 32'h85CFF0EF;
    mem['h0A96] <= 32'h00900613;
    mem['h0A97] <= 32'h01500593;
    mem['h0A98] <= 32'h01900513;
    mem['h0A99] <= 32'h84CFF0EF;
    mem['h0A9A] <= 32'hFDC42703;
    mem['h0A9B] <= 32'h00100793;
    mem['h0A9C] <= 32'h02F71A63;
    mem['h0A9D] <= 32'h00300613;
    mem['h0A9E] <= 32'h01500593;
    mem['h0A9F] <= 32'h00500513;
    mem['h0AA0] <= 32'h830FF0EF;
    mem['h0AA1] <= 32'h00900613;
    mem['h0AA2] <= 32'h01500593;
    mem['h0AA3] <= 32'h00F00513;
    mem['h0AA4] <= 32'h820FF0EF;
    mem['h0AA5] <= 32'h00900613;
    mem['h0AA6] <= 32'h01500593;
    mem['h0AA7] <= 32'h01900513;
    mem['h0AA8] <= 32'h810FF0EF;
    mem['h0AA9] <= 32'h00000013;
    mem['h0AAA] <= 32'h02C12083;
    mem['h0AAB] <= 32'h02812403;
    mem['h0AAC] <= 32'h03010113;
    mem['h0AAD] <= 32'h00008067;
    mem['h0AAE] <= 32'hFE010113;
    mem['h0AAF] <= 32'h00812E23;
    mem['h0AB0] <= 32'h02010413;
    mem['h0AB1] <= 32'h00800793;
    mem['h0AB2] <= 32'hFEF406A3;
    mem['h0AB3] <= 32'hFE0407A3;
    mem['h0AB4] <= 32'h4B00006F;
    mem['h0AB5] <= 32'hFE040723;
    mem['h0AB6] <= 32'h4900006F;
    mem['h0AB7] <= 32'hFEF44703;
    mem['h0AB8] <= 32'h00070793;
    mem['h0AB9] <= 32'h00279793;
    mem['h0ABA] <= 32'h00E787B3;
    mem['h0ABB] <= 32'h00379793;
    mem['h0ABC] <= 32'h00078713;
    mem['h0ABD] <= 32'hFEE44783;
    mem['h0ABE] <= 32'h00F707B3;
    mem['h0ABF] <= 32'h00279713;
    mem['h0AC0] <= 32'h052007B7;
    mem['h0AC1] <= 32'h00F707B3;
    mem['h0AC2] <= 32'h0007A023;
    mem['h0AC3] <= 32'hFEF44703;
    mem['h0AC4] <= 32'hFED44783;
    mem['h0AC5] <= 32'h00F71E63;
    mem['h0AC6] <= 32'hFEE44703;
    mem['h0AC7] <= 32'h00400793;
    mem['h0AC8] <= 32'h00E7F863;
    mem['h0AC9] <= 32'hFEE44703;
    mem['h0ACA] <= 32'h00700793;
    mem['h0ACB] <= 32'h02E7F663;
    mem['h0ACC] <= 32'hFEE44703;
    mem['h0ACD] <= 32'h00600793;
    mem['h0ACE] <= 32'h04F71A63;
    mem['h0ACF] <= 32'hFEF44703;
    mem['h0AD0] <= 32'hFED44783;
    mem['h0AD1] <= 32'h04F76463;
    mem['h0AD2] <= 32'hFEF44703;
    mem['h0AD3] <= 32'hFED44783;
    mem['h0AD4] <= 32'h00478793;
    mem['h0AD5] <= 32'h02E7CC63;
    mem['h0AD6] <= 32'hFEF44703;
    mem['h0AD7] <= 32'h00070793;
    mem['h0AD8] <= 32'h00279793;
    mem['h0AD9] <= 32'h00E787B3;
    mem['h0ADA] <= 32'h00379793;
    mem['h0ADB] <= 32'h00078713;
    mem['h0ADC] <= 32'hFEE44783;
    mem['h0ADD] <= 32'h00F707B3;
    mem['h0ADE] <= 32'h00279713;
    mem['h0ADF] <= 32'h052007B7;
    mem['h0AE0] <= 32'h00F707B3;
    mem['h0AE1] <= 32'h00300713;
    mem['h0AE2] <= 32'h00E7A023;
    mem['h0AE3] <= 32'hFEF44703;
    mem['h0AE4] <= 32'hFED44783;
    mem['h0AE5] <= 32'h00278793;
    mem['h0AE6] <= 32'h00F71E63;
    mem['h0AE7] <= 32'hFEE44703;
    mem['h0AE8] <= 32'h00800793;
    mem['h0AE9] <= 32'h00E7F863;
    mem['h0AEA] <= 32'hFEE44703;
    mem['h0AEB] <= 32'h00B00793;
    mem['h0AEC] <= 32'h02E7FC63;
    mem['h0AED] <= 32'hFEE44703;
    mem['h0AEE] <= 32'h00900793;
    mem['h0AEF] <= 32'h00F70863;
    mem['h0AF0] <= 32'hFEE44703;
    mem['h0AF1] <= 32'h00B00793;
    mem['h0AF2] <= 32'h04F71A63;
    mem['h0AF3] <= 32'hFEF44703;
    mem['h0AF4] <= 32'hFED44783;
    mem['h0AF5] <= 32'h04F76463;
    mem['h0AF6] <= 32'hFEF44703;
    mem['h0AF7] <= 32'hFED44783;
    mem['h0AF8] <= 32'h00478793;
    mem['h0AF9] <= 32'h02E7CC63;
    mem['h0AFA] <= 32'hFEF44703;
    mem['h0AFB] <= 32'h00070793;
    mem['h0AFC] <= 32'h00279793;
    mem['h0AFD] <= 32'h00E787B3;
    mem['h0AFE] <= 32'h00379793;
    mem['h0AFF] <= 32'h00078713;
    mem['h0B00] <= 32'hFEE44783;
    mem['h0B01] <= 32'h00F707B3;
    mem['h0B02] <= 32'h00279713;
    mem['h0B03] <= 32'h052007B7;
    mem['h0B04] <= 32'h00F707B3;
    mem['h0B05] <= 32'h00300713;
    mem['h0B06] <= 32'h00E7A023;
    mem['h0B07] <= 32'hFEF44703;
    mem['h0B08] <= 32'hFED44783;
    mem['h0B09] <= 32'h00F70A63;
    mem['h0B0A] <= 32'hFEF44703;
    mem['h0B0B] <= 32'hFED44783;
    mem['h0B0C] <= 32'h00478793;
    mem['h0B0D] <= 32'h00F71E63;
    mem['h0B0E] <= 32'hFEE44703;
    mem['h0B0F] <= 32'h00C00793;
    mem['h0B10] <= 32'h00E7F863;
    mem['h0B11] <= 32'hFEE44703;
    mem['h0B12] <= 32'h00F00793;
    mem['h0B13] <= 32'h04E7FA63;
    mem['h0B14] <= 32'hFEE44703;
    mem['h0B15] <= 32'h00D00793;
    mem['h0B16] <= 32'h02F71063;
    mem['h0B17] <= 32'hFEF44703;
    mem['h0B18] <= 32'hFED44783;
    mem['h0B19] <= 32'h00F76A63;
    mem['h0B1A] <= 32'hFEF44703;
    mem['h0B1B] <= 32'hFED44783;
    mem['h0B1C] <= 32'h00478793;
    mem['h0B1D] <= 32'h02E7D663;
    mem['h0B1E] <= 32'hFEF44703;
    mem['h0B1F] <= 32'hFED44783;
    mem['h0B20] <= 32'h00278793;
    mem['h0B21] <= 32'h04F71863;
    mem['h0B22] <= 32'hFEE44703;
    mem['h0B23] <= 32'h00C00793;
    mem['h0B24] <= 32'h04E7F263;
    mem['h0B25] <= 32'hFEE44703;
    mem['h0B26] <= 32'h00E00793;
    mem['h0B27] <= 32'h02E7EC63;
    mem['h0B28] <= 32'hFEF44703;
    mem['h0B29] <= 32'h00070793;
    mem['h0B2A] <= 32'h00279793;
    mem['h0B2B] <= 32'h00E787B3;
    mem['h0B2C] <= 32'h00379793;
    mem['h0B2D] <= 32'h00078713;
    mem['h0B2E] <= 32'hFEE44783;
    mem['h0B2F] <= 32'h00F707B3;
    mem['h0B30] <= 32'h00279713;
    mem['h0B31] <= 32'h052007B7;
    mem['h0B32] <= 32'h00F707B3;
    mem['h0B33] <= 32'h00300713;
    mem['h0B34] <= 32'h00E7A023;
    mem['h0B35] <= 32'hFEF44703;
    mem['h0B36] <= 32'hFED44783;
    mem['h0B37] <= 32'h00F70A63;
    mem['h0B38] <= 32'hFEF44703;
    mem['h0B39] <= 32'hFED44783;
    mem['h0B3A] <= 32'h00478793;
    mem['h0B3B] <= 32'h00F71E63;
    mem['h0B3C] <= 32'hFEE44703;
    mem['h0B3D] <= 32'h01300793;
    mem['h0B3E] <= 32'h00E7F863;
    mem['h0B3F] <= 32'hFEE44703;
    mem['h0B40] <= 32'h01600793;
    mem['h0B41] <= 32'h04E7FA63;
    mem['h0B42] <= 32'hFEE44703;
    mem['h0B43] <= 32'h01400793;
    mem['h0B44] <= 32'h02F71063;
    mem['h0B45] <= 32'hFEF44703;
    mem['h0B46] <= 32'hFED44783;
    mem['h0B47] <= 32'h00F76A63;
    mem['h0B48] <= 32'hFEF44703;
    mem['h0B49] <= 32'hFED44783;
    mem['h0B4A] <= 32'h00478793;
    mem['h0B4B] <= 32'h02E7D663;
    mem['h0B4C] <= 32'hFEF44703;
    mem['h0B4D] <= 32'hFED44783;
    mem['h0B4E] <= 32'h00278793;
    mem['h0B4F] <= 32'h04F71863;
    mem['h0B50] <= 32'hFEE44703;
    mem['h0B51] <= 32'h01300793;
    mem['h0B52] <= 32'h04E7F263;
    mem['h0B53] <= 32'hFEE44703;
    mem['h0B54] <= 32'h01500793;
    mem['h0B55] <= 32'h02E7EC63;
    mem['h0B56] <= 32'hFEF44703;
    mem['h0B57] <= 32'h00070793;
    mem['h0B58] <= 32'h00279793;
    mem['h0B59] <= 32'h00E787B3;
    mem['h0B5A] <= 32'h00379793;
    mem['h0B5B] <= 32'h00078713;
    mem['h0B5C] <= 32'hFEE44783;
    mem['h0B5D] <= 32'h00F707B3;
    mem['h0B5E] <= 32'h00279713;
    mem['h0B5F] <= 32'h052007B7;
    mem['h0B60] <= 32'h00F707B3;
    mem['h0B61] <= 32'h00300713;
    mem['h0B62] <= 32'h00E7A023;
    mem['h0B63] <= 32'hFEF44703;
    mem['h0B64] <= 32'hFED44783;
    mem['h0B65] <= 32'h00278793;
    mem['h0B66] <= 32'h00F71863;
    mem['h0B67] <= 32'hFEE44703;
    mem['h0B68] <= 32'h01900793;
    mem['h0B69] <= 32'h04F70A63;
    mem['h0B6A] <= 32'hFEF44703;
    mem['h0B6B] <= 32'hFED44783;
    mem['h0B6C] <= 32'h00378793;
    mem['h0B6D] <= 32'h00F71863;
    mem['h0B6E] <= 32'hFEE44703;
    mem['h0B6F] <= 32'h01A00793;
    mem['h0B70] <= 32'h02F70C63;
    mem['h0B71] <= 32'hFEE44703;
    mem['h0B72] <= 32'h01800793;
    mem['h0B73] <= 32'h00F70863;
    mem['h0B74] <= 32'hFEE44703;
    mem['h0B75] <= 32'h01B00793;
    mem['h0B76] <= 32'h04F71A63;
    mem['h0B77] <= 32'hFEF44703;
    mem['h0B78] <= 32'hFED44783;
    mem['h0B79] <= 32'h04F76463;
    mem['h0B7A] <= 32'hFEF44703;
    mem['h0B7B] <= 32'hFED44783;
    mem['h0B7C] <= 32'h00478793;
    mem['h0B7D] <= 32'h02E7CC63;
    mem['h0B7E] <= 32'hFEF44703;
    mem['h0B7F] <= 32'h00070793;
    mem['h0B80] <= 32'h00279793;
    mem['h0B81] <= 32'h00E787B3;
    mem['h0B82] <= 32'h00379793;
    mem['h0B83] <= 32'h00078713;
    mem['h0B84] <= 32'hFEE44783;
    mem['h0B85] <= 32'h00F707B3;
    mem['h0B86] <= 32'h00279713;
    mem['h0B87] <= 32'h052007B7;
    mem['h0B88] <= 32'h00F707B3;
    mem['h0B89] <= 32'h00300713;
    mem['h0B8A] <= 32'h00E7A023;
    mem['h0B8B] <= 32'hFEE44703;
    mem['h0B8C] <= 32'h01F00793;
    mem['h0B8D] <= 32'h02F71063;
    mem['h0B8E] <= 32'hFED44703;
    mem['h0B8F] <= 32'hFEF44783;
    mem['h0B90] <= 32'h00F77A63;
    mem['h0B91] <= 32'hFEF44703;
    mem['h0B92] <= 32'hFED44783;
    mem['h0B93] <= 32'h00378793;
    mem['h0B94] <= 32'h06E7D063;
    mem['h0B95] <= 32'hFEF44703;
    mem['h0B96] <= 32'hFED44783;
    mem['h0B97] <= 32'h00F70A63;
    mem['h0B98] <= 32'hFEF44703;
    mem['h0B99] <= 32'hFED44783;
    mem['h0B9A] <= 32'h00478793;
    mem['h0B9B] <= 32'h00F71E63;
    mem['h0B9C] <= 32'hFEE44703;
    mem['h0B9D] <= 32'h01C00793;
    mem['h0B9E] <= 32'h00E7F863;
    mem['h0B9F] <= 32'hFEE44703;
    mem['h0BA0] <= 32'h01E00793;
    mem['h0BA1] <= 32'h02E7F663;
    mem['h0BA2] <= 32'hFEE44703;
    mem['h0BA3] <= 32'h01D00793;
    mem['h0BA4] <= 32'h04F71A63;
    mem['h0BA5] <= 32'hFEF44703;
    mem['h0BA6] <= 32'hFED44783;
    mem['h0BA7] <= 32'h04F76463;
    mem['h0BA8] <= 32'hFEF44703;
    mem['h0BA9] <= 32'hFED44783;
    mem['h0BAA] <= 32'h00478793;
    mem['h0BAB] <= 32'h02E7CC63;
    mem['h0BAC] <= 32'hFEF44703;
    mem['h0BAD] <= 32'h00070793;
    mem['h0BAE] <= 32'h00279793;
    mem['h0BAF] <= 32'h00E787B3;
    mem['h0BB0] <= 32'h00379793;
    mem['h0BB1] <= 32'h00078713;
    mem['h0BB2] <= 32'hFEE44783;
    mem['h0BB3] <= 32'h00F707B3;
    mem['h0BB4] <= 32'h00279713;
    mem['h0BB5] <= 32'h052007B7;
    mem['h0BB6] <= 32'h00F707B3;
    mem['h0BB7] <= 32'h00300713;
    mem['h0BB8] <= 32'h00E7A023;
    mem['h0BB9] <= 32'hFEE44703;
    mem['h0BBA] <= 32'h02100793;
    mem['h0BBB] <= 32'h02F71063;
    mem['h0BBC] <= 32'hFEF44703;
    mem['h0BBD] <= 32'hFED44783;
    mem['h0BBE] <= 32'h00F76A63;
    mem['h0BBF] <= 32'hFEF44703;
    mem['h0BC0] <= 32'hFED44783;
    mem['h0BC1] <= 32'h00278793;
    mem['h0BC2] <= 32'h02E7D063;
    mem['h0BC3] <= 32'hFEE44703;
    mem['h0BC4] <= 32'h02100793;
    mem['h0BC5] <= 32'h04F71463;
    mem['h0BC6] <= 32'hFEF44703;
    mem['h0BC7] <= 32'hFED44783;
    mem['h0BC8] <= 32'h00478793;
    mem['h0BC9] <= 32'h02F71C63;
    mem['h0BCA] <= 32'hFEF44703;
    mem['h0BCB] <= 32'h00070793;
    mem['h0BCC] <= 32'h00279793;
    mem['h0BCD] <= 32'h00E787B3;
    mem['h0BCE] <= 32'h00379793;
    mem['h0BCF] <= 32'h00078713;
    mem['h0BD0] <= 32'hFEE44783;
    mem['h0BD1] <= 32'h00F707B3;
    mem['h0BD2] <= 32'h00279713;
    mem['h0BD3] <= 32'h052007B7;
    mem['h0BD4] <= 32'h00F707B3;
    mem['h0BD5] <= 32'h00300713;
    mem['h0BD6] <= 32'h00E7A023;
    mem['h0BD7] <= 32'hFEE44783;
    mem['h0BD8] <= 32'h00178793;
    mem['h0BD9] <= 32'hFEF40723;
    mem['h0BDA] <= 32'hFEE44703;
    mem['h0BDB] <= 32'h02700793;
    mem['h0BDC] <= 32'hB6E7F6E3;
    mem['h0BDD] <= 32'hFEF44783;
    mem['h0BDE] <= 32'h00178793;
    mem['h0BDF] <= 32'hFEF407A3;
    mem['h0BE0] <= 32'hFEF44703;
    mem['h0BE1] <= 32'h01600793;
    mem['h0BE2] <= 32'hB4E7F6E3;
    mem['h0BE3] <= 32'h00000013;
    mem['h0BE4] <= 32'h00000013;
    mem['h0BE5] <= 32'h01C12403;
    mem['h0BE6] <= 32'h02010113;
    mem['h0BE7] <= 32'h00008067;
    mem['h0BE8] <= 32'hFE010113;
    mem['h0BE9] <= 32'h00812E23;
    mem['h0BEA] <= 32'h02010413;
    mem['h0BEB] <= 32'h000017B7;
    mem['h0BEC] <= 32'hFFF78793;
    mem['h0BED] <= 32'hFEF42623;
    mem['h0BEE] <= 32'hFE0405A3;
    mem['h0BEF] <= 32'h4D40006F;
    mem['h0BF0] <= 32'hFE040523;
    mem['h0BF1] <= 32'h4B40006F;
    mem['h0BF2] <= 32'hFE0404A3;
    mem['h0BF3] <= 32'h4940006F;
    mem['h0BF4] <= 32'hFEB44783;
    mem['h0BF5] <= 32'h04079863;
    mem['h0BF6] <= 32'hFEA44783;
    mem['h0BF7] <= 32'h00078863;
    mem['h0BF8] <= 32'hFEA44703;
    mem['h0BF9] <= 32'h00100793;
    mem['h0BFA] <= 32'h00F71863;
    mem['h0BFB] <= 32'h22200793;
    mem['h0BFC] <= 32'hFEF42623;
    mem['h0BFD] <= 32'h4300006F;
    mem['h0BFE] <= 32'hFE944703;
    mem['h0BFF] <= 32'h00E00793;
    mem['h0C00] <= 32'h00F70863;
    mem['h0C01] <= 32'hFE944703;
    mem['h0C02] <= 32'h00F00793;
    mem['h0C03] <= 32'h00F71863;
    mem['h0C04] <= 32'h11100793;
    mem['h0C05] <= 32'hFEF42623;
    mem['h0C06] <= 32'h40C0006F;
    mem['h0C07] <= 32'hFE042623;
    mem['h0C08] <= 32'h4040006F;
    mem['h0C09] <= 32'hFEB44703;
    mem['h0C0A] <= 32'h00100793;
    mem['h0C0B] <= 32'h04F71C63;
    mem['h0C0C] <= 32'hFEA44783;
    mem['h0C0D] <= 32'h00078863;
    mem['h0C0E] <= 32'hFEA44703;
    mem['h0C0F] <= 32'h00100793;
    mem['h0C10] <= 32'h00F71863;
    mem['h0C11] <= 32'h08000793;
    mem['h0C12] <= 32'hFEF42623;
    mem['h0C13] <= 32'h3D80006F;
    mem['h0C14] <= 32'hFE944703;
    mem['h0C15] <= 32'h00E00793;
    mem['h0C16] <= 32'h00F70863;
    mem['h0C17] <= 32'hFE944703;
    mem['h0C18] <= 32'h00F00793;
    mem['h0C19] <= 32'h00F71863;
    mem['h0C1A] <= 32'h08000793;
    mem['h0C1B] <= 32'hFEF42623;
    mem['h0C1C] <= 32'h3B40006F;
    mem['h0C1D] <= 32'h000017B7;
    mem['h0C1E] <= 32'h8B478793;
    mem['h0C1F] <= 32'hFEF42623;
    mem['h0C20] <= 32'h3A40006F;
    mem['h0C21] <= 32'hFEB44703;
    mem['h0C22] <= 32'h00200793;
    mem['h0C23] <= 32'h04F71A63;
    mem['h0C24] <= 32'hFEA44783;
    mem['h0C25] <= 32'h00078863;
    mem['h0C26] <= 32'hFEA44703;
    mem['h0C27] <= 32'h00100793;
    mem['h0C28] <= 32'h00F71863;
    mem['h0C29] <= 32'h00B00793;
    mem['h0C2A] <= 32'hFEF42623;
    mem['h0C2B] <= 32'h3780006F;
    mem['h0C2C] <= 32'hFE944703;
    mem['h0C2D] <= 32'h00E00793;
    mem['h0C2E] <= 32'h00F70863;
    mem['h0C2F] <= 32'hFE944703;
    mem['h0C30] <= 32'h00F00793;
    mem['h0C31] <= 32'h00F71863;
    mem['h0C32] <= 32'h00B00793;
    mem['h0C33] <= 32'hFEF42623;
    mem['h0C34] <= 32'h3540006F;
    mem['h0C35] <= 32'h00900793;
    mem['h0C36] <= 32'hFEF42623;
    mem['h0C37] <= 32'h3480006F;
    mem['h0C38] <= 32'hFEB44703;
    mem['h0C39] <= 32'h00300793;
    mem['h0C3A] <= 32'h06F71063;
    mem['h0C3B] <= 32'hFEA44783;
    mem['h0C3C] <= 32'h00078863;
    mem['h0C3D] <= 32'hFEA44703;
    mem['h0C3E] <= 32'h00100793;
    mem['h0C3F] <= 32'h00F71A63;
    mem['h0C40] <= 32'h000017B7;
    mem['h0C41] <= 32'hA0078793;
    mem['h0C42] <= 32'hFEF42623;
    mem['h0C43] <= 32'h3180006F;
    mem['h0C44] <= 32'hFE944703;
    mem['h0C45] <= 32'h00E00793;
    mem['h0C46] <= 32'h00F70863;
    mem['h0C47] <= 32'hFE944703;
    mem['h0C48] <= 32'h00F00793;
    mem['h0C49] <= 32'h00F71A63;
    mem['h0C4A] <= 32'h000017B7;
    mem['h0C4B] <= 32'hB0078793;
    mem['h0C4C] <= 32'hFEF42623;
    mem['h0C4D] <= 32'h2F00006F;
    mem['h0C4E] <= 32'h000017B7;
    mem['h0C4F] <= 32'hF0078793;
    mem['h0C50] <= 32'hFEF42623;
    mem['h0C51] <= 32'h2E00006F;
    mem['h0C52] <= 32'hFEB44703;
    mem['h0C53] <= 32'h00400793;
    mem['h0C54] <= 32'h06F71063;
    mem['h0C55] <= 32'hFEA44783;
    mem['h0C56] <= 32'h00078863;
    mem['h0C57] <= 32'hFEA44703;
    mem['h0C58] <= 32'h00100793;
    mem['h0C59] <= 32'h00F71A63;
    mem['h0C5A] <= 32'h000017B7;
    mem['h0C5B] <= 32'hFD878793;
    mem['h0C5C] <= 32'hFEF42623;
    mem['h0C5D] <= 32'h2B00006F;
    mem['h0C5E] <= 32'hFE944703;
    mem['h0C5F] <= 32'h00E00793;
    mem['h0C60] <= 32'h00F70863;
    mem['h0C61] <= 32'hFE944703;
    mem['h0C62] <= 32'h00F00793;
    mem['h0C63] <= 32'h00F71A63;
    mem['h0C64] <= 32'h000017B7;
    mem['h0C65] <= 32'hFD478793;
    mem['h0C66] <= 32'hFEF42623;
    mem['h0C67] <= 32'h2880006F;
    mem['h0C68] <= 32'h000017B7;
    mem['h0C69] <= 32'hFF078793;
    mem['h0C6A] <= 32'hFEF42623;
    mem['h0C6B] <= 32'h2780006F;
    mem['h0C6C] <= 32'hFEB44703;
    mem['h0C6D] <= 32'h00500793;
    mem['h0C6E] <= 32'h04F71A63;
    mem['h0C6F] <= 32'hFEA44783;
    mem['h0C70] <= 32'h00078863;
    mem['h0C71] <= 32'hFEA44703;
    mem['h0C72] <= 32'h00100793;
    mem['h0C73] <= 32'h00F71863;
    mem['h0C74] <= 32'h75D00793;
    mem['h0C75] <= 32'hFEF42623;
    mem['h0C76] <= 32'h24C0006F;
    mem['h0C77] <= 32'hFE944703;
    mem['h0C78] <= 32'h00E00793;
    mem['h0C79] <= 32'h00F70863;
    mem['h0C7A] <= 32'hFE944703;
    mem['h0C7B] <= 32'h00F00793;
    mem['h0C7C] <= 32'h00F71863;
    mem['h0C7D] <= 32'h74D00793;
    mem['h0C7E] <= 32'hFEF42623;
    mem['h0C7F] <= 32'h2280006F;
    mem['h0C80] <= 32'h70D00793;
    mem['h0C81] <= 32'hFEF42623;
    mem['h0C82] <= 32'h21C0006F;
    mem['h0C83] <= 32'hFEB44703;
    mem['h0C84] <= 32'h00600793;
    mem['h0C85] <= 32'h06F71063;
    mem['h0C86] <= 32'hFEA44783;
    mem['h0C87] <= 32'h00078863;
    mem['h0C88] <= 32'hFEA44703;
    mem['h0C89] <= 32'h00100793;
    mem['h0C8A] <= 32'h00F71A63;
    mem['h0C8B] <= 32'h000017B7;
    mem['h0C8C] <= 32'hFAF78793;
    mem['h0C8D] <= 32'hFEF42623;
    mem['h0C8E] <= 32'h1EC0006F;
    mem['h0C8F] <= 32'hFE944703;
    mem['h0C90] <= 32'h00E00793;
    mem['h0C91] <= 32'h00F70863;
    mem['h0C92] <= 32'hFE944703;
    mem['h0C93] <= 32'h00F00793;
    mem['h0C94] <= 32'h00F71A63;
    mem['h0C95] <= 32'h000017B7;
    mem['h0C96] <= 32'hF6F78793;
    mem['h0C97] <= 32'hFEF42623;
    mem['h0C98] <= 32'h1C40006F;
    mem['h0C99] <= 32'h000017B7;
    mem['h0C9A] <= 32'hF0F78793;
    mem['h0C9B] <= 32'hFEF42623;
    mem['h0C9C] <= 32'h1B40006F;
    mem['h0C9D] <= 32'hFEB44703;
    mem['h0C9E] <= 32'h00700793;
    mem['h0C9F] <= 32'h06F71063;
    mem['h0CA0] <= 32'hFEA44783;
    mem['h0CA1] <= 32'h00078863;
    mem['h0CA2] <= 32'hFEA44703;
    mem['h0CA3] <= 32'h00100793;
    mem['h0CA4] <= 32'h00F71A63;
    mem['h0CA5] <= 32'h000017B7;
    mem['h0CA6] <= 32'hFB078793;
    mem['h0CA7] <= 32'hFEF42623;
    mem['h0CA8] <= 32'h1840006F;
    mem['h0CA9] <= 32'hFE944703;
    mem['h0CAA] <= 32'h00E00793;
    mem['h0CAB] <= 32'h00F70863;
    mem['h0CAC] <= 32'hFE944703;
    mem['h0CAD] <= 32'h00F00793;
    mem['h0CAE] <= 32'h00F71A63;
    mem['h0CAF] <= 32'h000017B7;
    mem['h0CB0] <= 32'hF9078793;
    mem['h0CB1] <= 32'hFEF42623;
    mem['h0CB2] <= 32'h15C0006F;
    mem['h0CB3] <= 32'h000017B7;
    mem['h0CB4] <= 32'hFA078793;
    mem['h0CB5] <= 32'hFEF42623;
    mem['h0CB6] <= 32'h14C0006F;
    mem['h0CB7] <= 32'hFEB44703;
    mem['h0CB8] <= 32'h00800793;
    mem['h0CB9] <= 32'h00F71863;
    mem['h0CBA] <= 32'h0A000793;
    mem['h0CBB] <= 32'hFEF42623;
    mem['h0CBC] <= 32'h1340006F;
    mem['h0CBD] <= 32'hFEB44703;
    mem['h0CBE] <= 32'h00900793;
    mem['h0CBF] <= 32'h04F71E63;
    mem['h0CC0] <= 32'hFE944703;
    mem['h0CC1] <= 32'h00E00793;
    mem['h0CC2] <= 32'h00F70863;
    mem['h0CC3] <= 32'hFE944703;
    mem['h0CC4] <= 32'h00F00793;
    mem['h0CC5] <= 32'h00F71A63;
    mem['h0CC6] <= 32'h000017B7;
    mem['h0CC7] <= 32'hCCC78793;
    mem['h0CC8] <= 32'hFEF42623;
    mem['h0CC9] <= 32'h1000006F;
    mem['h0CCA] <= 32'hFEA44783;
    mem['h0CCB] <= 32'h00078863;
    mem['h0CCC] <= 32'hFEA44703;
    mem['h0CCD] <= 32'h00100793;
    mem['h0CCE] <= 32'h00F71863;
    mem['h0CCF] <= 32'h11100793;
    mem['h0CD0] <= 32'hFEF42623;
    mem['h0CD1] <= 32'h0E00006F;
    mem['h0CD2] <= 32'h000017B7;
    mem['h0CD3] <= 32'hAAA78793;
    mem['h0CD4] <= 32'hFEF42623;
    mem['h0CD5] <= 32'h0D00006F;
    mem['h0CD6] <= 32'hFEB44703;
    mem['h0CD7] <= 32'h00A00793;
    mem['h0CD8] <= 32'h04F71A63;
    mem['h0CD9] <= 32'hFEA44783;
    mem['h0CDA] <= 32'h00078863;
    mem['h0CDB] <= 32'hFEA44703;
    mem['h0CDC] <= 32'h00100793;
    mem['h0CDD] <= 32'h00F71863;
    mem['h0CDE] <= 32'h00B00793;
    mem['h0CDF] <= 32'hFEF42623;
    mem['h0CE0] <= 32'h0A40006F;
    mem['h0CE1] <= 32'hFE944703;
    mem['h0CE2] <= 32'h00E00793;
    mem['h0CE3] <= 32'h00F70863;
    mem['h0CE4] <= 32'hFE944703;
    mem['h0CE5] <= 32'h00F00793;
    mem['h0CE6] <= 32'h00F71863;
    mem['h0CE7] <= 32'h00B00793;
    mem['h0CE8] <= 32'hFEF42623;
    mem['h0CE9] <= 32'h0800006F;
    mem['h0CEA] <= 32'h00700793;
    mem['h0CEB] <= 32'hFEF42623;
    mem['h0CEC] <= 32'h0740006F;
    mem['h0CED] <= 32'hFEB44703;
    mem['h0CEE] <= 32'h00B00793;
    mem['h0CEF] <= 32'h00F71A63;
    mem['h0CF0] <= 32'h000017B7;
    mem['h0CF1] <= 32'hAA078793;
    mem['h0CF2] <= 32'hFEF42623;
    mem['h0CF3] <= 32'h0580006F;
    mem['h0CF4] <= 32'hFEB44703;
    mem['h0CF5] <= 32'h00C00793;
    mem['h0CF6] <= 32'h00F71863;
    mem['h0CF7] <= 32'h0AA00793;
    mem['h0CF8] <= 32'hFEF42623;
    mem['h0CF9] <= 32'h0400006F;
    mem['h0CFA] <= 32'hFEB44703;
    mem['h0CFB] <= 32'h00D00793;
    mem['h0CFC] <= 32'h00F71A63;
    mem['h0CFD] <= 32'h000017B7;
    mem['h0CFE] <= 32'hA0A78793;
    mem['h0CFF] <= 32'hFEF42623;
    mem['h0D00] <= 32'h0240006F;
    mem['h0D01] <= 32'hFEB44703;
    mem['h0D02] <= 32'h00E00793;
    mem['h0D03] <= 32'h00F71A63;
    mem['h0D04] <= 32'h000017B7;
    mem['h0D05] <= 32'hFFF78793;
    mem['h0D06] <= 32'hFEF42623;
    mem['h0D07] <= 32'h0080006F;
    mem['h0D08] <= 32'hFE042623;
    mem['h0D09] <= 32'hFEB44783;
    mem['h0D0A] <= 32'h00479713;
    mem['h0D0B] <= 32'hFEA44783;
    mem['h0D0C] <= 32'h00F707B3;
    mem['h0D0D] <= 32'h00479713;
    mem['h0D0E] <= 32'hFE944783;
    mem['h0D0F] <= 32'h00F707B3;
    mem['h0D10] <= 32'h00279713;
    mem['h0D11] <= 32'h051007B7;
    mem['h0D12] <= 32'h00F707B3;
    mem['h0D13] <= 32'hFEC42703;
    mem['h0D14] <= 32'h00E7A023;
    mem['h0D15] <= 32'hFE944783;
    mem['h0D16] <= 32'h00178793;
    mem['h0D17] <= 32'hFEF404A3;
    mem['h0D18] <= 32'hFE944703;
    mem['h0D19] <= 32'h00F00793;
    mem['h0D1A] <= 32'hB6E7F4E3;
    mem['h0D1B] <= 32'hFEA44783;
    mem['h0D1C] <= 32'h00178793;
    mem['h0D1D] <= 32'hFEF40523;
    mem['h0D1E] <= 32'hFEA44703;
    mem['h0D1F] <= 32'h00F00793;
    mem['h0D20] <= 32'hB4E7F4E3;
    mem['h0D21] <= 32'hFEB44783;
    mem['h0D22] <= 32'h00178793;
    mem['h0D23] <= 32'hFEF405A3;
    mem['h0D24] <= 32'hFEB44703;
    mem['h0D25] <= 32'h00F00793;
    mem['h0D26] <= 32'hB2E7F4E3;
    mem['h0D27] <= 32'h00000013;
    mem['h0D28] <= 32'h00000013;
    mem['h0D29] <= 32'h01C12403;
    mem['h0D2A] <= 32'h02010113;
    mem['h0D2B] <= 32'h00008067;
    mem['h0D2C] <= 32'hFD010113;
    mem['h0D2D] <= 32'h02812623;
    mem['h0D2E] <= 32'h03010413;
    mem['h0D2F] <= 32'hFCA42E23;
    mem['h0D30] <= 32'hFCB42C23;
    mem['h0D31] <= 32'hFCC42A23;
    mem['h0D32] <= 32'hFE042623;
    mem['h0D33] <= 32'hFD442703;
    mem['h0D34] <= 32'h41F75793;
    mem['h0D35] <= 32'h01E7D793;
    mem['h0D36] <= 32'h00F70733;
    mem['h0D37] <= 32'h00377713;
    mem['h0D38] <= 32'h40F707B3;
    mem['h0D39] <= 32'h00300713;
    mem['h0D3A] <= 32'h08E78063;
    mem['h0D3B] <= 32'h00300713;
    mem['h0D3C] <= 32'h08F74C63;
    mem['h0D3D] <= 32'h00200713;
    mem['h0D3E] <= 32'h04E78863;
    mem['h0D3F] <= 32'h00200713;
    mem['h0D40] <= 32'h08F74463;
    mem['h0D41] <= 32'h00078863;
    mem['h0D42] <= 32'h00100713;
    mem['h0D43] <= 32'h02E78063;
    mem['h0D44] <= 32'h0780006F;
    mem['h0D45] <= 32'hFD842783;
    mem['h0D46] <= 32'h00279793;
    mem['h0D47] <= 32'hFDC42703;
    mem['h0D48] <= 32'h00F707B3;
    mem['h0D49] <= 32'hFEF42623;
    mem['h0D4A] <= 32'h0600006F;
    mem['h0D4B] <= 32'hFD842783;
    mem['h0D4C] <= 32'h00C78713;
    mem['h0D4D] <= 32'hFDC42783;
    mem['h0D4E] <= 32'h00279793;
    mem['h0D4F] <= 32'h40F707B3;
    mem['h0D50] <= 32'hFEF42623;
    mem['h0D51] <= 32'h0440006F;
    mem['h0D52] <= 32'hFD842783;
    mem['h0D53] <= 32'h00279793;
    mem['h0D54] <= 32'h00F00713;
    mem['h0D55] <= 32'h40F70733;
    mem['h0D56] <= 32'hFDC42783;
    mem['h0D57] <= 32'h40F707B3;
    mem['h0D58] <= 32'hFEF42623;
    mem['h0D59] <= 32'h0240006F;
    mem['h0D5A] <= 32'h00300713;
    mem['h0D5B] <= 32'hFD842783;
    mem['h0D5C] <= 32'h40F70733;
    mem['h0D5D] <= 32'hFDC42783;
    mem['h0D5E] <= 32'h00279793;
    mem['h0D5F] <= 32'h00F707B3;
    mem['h0D60] <= 32'hFEF42623;
    mem['h0D61] <= 32'h00000013;
    mem['h0D62] <= 32'hFEC42783;
    mem['h0D63] <= 32'h00078513;
    mem['h0D64] <= 32'h02C12403;
    mem['h0D65] <= 32'h03010113;
    mem['h0D66] <= 32'h00008067;
    mem['h0D67] <= 32'hFD010113;
    mem['h0D68] <= 32'h02112623;
    mem['h0D69] <= 32'h02812423;
    mem['h0D6A] <= 32'h03010413;
    mem['h0D6B] <= 32'hFCA42E23;
    mem['h0D6C] <= 32'hFCB42C23;
    mem['h0D6D] <= 32'hFCC42A23;
    mem['h0D6E] <= 32'hFCD42823;
    mem['h0D6F] <= 32'hFE042623;
    mem['h0D70] <= 32'h0FC0006F;
    mem['h0D71] <= 32'hFE042423;
    mem['h0D72] <= 32'h0DC0006F;
    mem['h0D73] <= 32'hFD842603;
    mem['h0D74] <= 32'hFE842583;
    mem['h0D75] <= 32'hFEC42503;
    mem['h0D76] <= 32'hED9FF0EF;
    mem['h0D77] <= 32'hFEA42223;
    mem['h0D78] <= 32'hFD042703;
    mem['h0D79] <= 32'hFE842783;
    mem['h0D7A] <= 32'h00F70733;
    mem['h0D7B] <= 32'h00070793;
    mem['h0D7C] <= 32'h00279793;
    mem['h0D7D] <= 32'h00E787B3;
    mem['h0D7E] <= 32'h00379793;
    mem['h0D7F] <= 32'h00078693;
    mem['h0D80] <= 32'hFD442703;
    mem['h0D81] <= 32'hFEC42783;
    mem['h0D82] <= 32'h00F707B3;
    mem['h0D83] <= 32'h00F687B3;
    mem['h0D84] <= 32'hFEF42023;
    mem['h0D85] <= 32'hFD442703;
    mem['h0D86] <= 32'hFEC42783;
    mem['h0D87] <= 32'h00F707B3;
    mem['h0D88] <= 32'h0607CC63;
    mem['h0D89] <= 32'hFD442703;
    mem['h0D8A] <= 32'hFEC42783;
    mem['h0D8B] <= 32'h00F70733;
    mem['h0D8C] <= 32'h02700793;
    mem['h0D8D] <= 32'h06E7C263;
    mem['h0D8E] <= 32'hFD042703;
    mem['h0D8F] <= 32'hFE842783;
    mem['h0D90] <= 32'h00F707B3;
    mem['h0D91] <= 32'h0407CA63;
    mem['h0D92] <= 32'hFD042703;
    mem['h0D93] <= 32'hFE842783;
    mem['h0D94] <= 32'h00F70733;
    mem['h0D95] <= 32'h01D00793;
    mem['h0D96] <= 32'h04E7C063;
    mem['h0D97] <= 32'h00000713;
    mem['h0D98] <= 32'hFDC42783;
    mem['h0D99] <= 32'h00479793;
    mem['h0D9A] <= 32'h00F70733;
    mem['h0D9B] <= 32'hFE442783;
    mem['h0D9C] <= 32'h00F707B3;
    mem['h0D9D] <= 32'h0007C783;
    mem['h0D9E] <= 32'h02078063;
    mem['h0D9F] <= 32'h07C00713;
    mem['h0DA0] <= 32'hFE042783;
    mem['h0DA1] <= 32'h00F707B3;
    mem['h0DA2] <= 32'h0007C783;
    mem['h0DA3] <= 32'h00078663;
    mem['h0DA4] <= 32'h00000793;
    mem['h0DA5] <= 32'h0380006F;
    mem['h0DA6] <= 32'hFE842783;
    mem['h0DA7] <= 32'h00178793;
    mem['h0DA8] <= 32'hFEF42423;
    mem['h0DA9] <= 32'hFE842703;
    mem['h0DAA] <= 32'h00300793;
    mem['h0DAB] <= 32'hF2E7D0E3;
    mem['h0DAC] <= 32'hFEC42783;
    mem['h0DAD] <= 32'h00178793;
    mem['h0DAE] <= 32'hFEF42623;
    mem['h0DAF] <= 32'hFEC42703;
    mem['h0DB0] <= 32'h00300793;
    mem['h0DB1] <= 32'hF0E7D0E3;
    mem['h0DB2] <= 32'h00100793;
    mem['h0DB3] <= 32'h00078513;
    mem['h0DB4] <= 32'h02C12083;
    mem['h0DB5] <= 32'h02812403;
    mem['h0DB6] <= 32'h03010113;
    mem['h0DB7] <= 32'h00008067;
    mem['h0DB8] <= 32'hFD010113;
    mem['h0DB9] <= 32'h02812623;
    mem['h0DBA] <= 32'h03010413;
    mem['h0DBB] <= 32'hFCA42E23;
    mem['h0DBC] <= 32'hFCB42C23;
    mem['h0DBD] <= 32'hFCC42A23;
    mem['h0DBE] <= 32'hFD442783;
    mem['h0DBF] <= 32'hFEF407A3;
    mem['h0DC0] <= 32'h7000006F;
    mem['h0DC1] <= 32'hFD842783;
    mem['h0DC2] <= 32'hFEF40723;
    mem['h0DC3] <= 32'h6D80006F;
    mem['h0DC4] <= 32'hFDC42703;
    mem['h0DC5] <= 32'h00900793;
    mem['h0DC6] <= 32'h6AE7EE63;
    mem['h0DC7] <= 32'hFDC42783;
    mem['h0DC8] <= 32'h00279713;
    mem['h0DC9] <= 32'h001057B7;
    mem['h0DCA] <= 32'h45C78793;
    mem['h0DCB] <= 32'h00F707B3;
    mem['h0DCC] <= 32'h0007A783;
    mem['h0DCD] <= 32'h00078067;
    mem['h0DCE] <= 32'hFEE44783;
    mem['h0DCF] <= 32'hFD842703;
    mem['h0DD0] <= 32'h02F70863;
    mem['h0DD1] <= 32'hFEE44703;
    mem['h0DD2] <= 32'hFD842783;
    mem['h0DD3] <= 32'h00278793;
    mem['h0DD4] <= 32'h02F70063;
    mem['h0DD5] <= 32'hFEF44783;
    mem['h0DD6] <= 32'hFD442703;
    mem['h0DD7] <= 32'h00F70A63;
    mem['h0DD8] <= 32'hFEF44703;
    mem['h0DD9] <= 32'hFD442783;
    mem['h0DDA] <= 32'h00478793;
    mem['h0DDB] <= 32'h02F71A63;
    mem['h0DDC] <= 32'hFEF44703;
    mem['h0DDD] <= 32'h00070793;
    mem['h0DDE] <= 32'h00279793;
    mem['h0DDF] <= 32'h00E787B3;
    mem['h0DE0] <= 32'h00379793;
    mem['h0DE1] <= 32'h00078713;
    mem['h0DE2] <= 32'hFEE44783;
    mem['h0DE3] <= 32'h00F707B3;
    mem['h0DE4] <= 32'h07C00713;
    mem['h0DE5] <= 32'h00F707B3;
    mem['h0DE6] <= 32'h00078023;
    mem['h0DE7] <= 32'h63C0006F;
    mem['h0DE8] <= 32'hFEF44703;
    mem['h0DE9] <= 32'h00070793;
    mem['h0DEA] <= 32'h00279793;
    mem['h0DEB] <= 32'h00E787B3;
    mem['h0DEC] <= 32'h00379793;
    mem['h0DED] <= 32'h00078713;
    mem['h0DEE] <= 32'hFEE44783;
    mem['h0DEF] <= 32'h00F707B3;
    mem['h0DF0] <= 32'h07C00713;
    mem['h0DF1] <= 32'h00F707B3;
    mem['h0DF2] <= 32'h00900713;
    mem['h0DF3] <= 32'h00E78023;
    mem['h0DF4] <= 32'h6080006F;
    mem['h0DF5] <= 32'hFEE44703;
    mem['h0DF6] <= 32'hFD842783;
    mem['h0DF7] <= 32'h00278793;
    mem['h0DF8] <= 32'h00F70A63;
    mem['h0DF9] <= 32'hFEF44703;
    mem['h0DFA] <= 32'hFD442783;
    mem['h0DFB] <= 32'h00178793;
    mem['h0DFC] <= 32'h02F71A63;
    mem['h0DFD] <= 32'hFEF44703;
    mem['h0DFE] <= 32'h00070793;
    mem['h0DFF] <= 32'h00279793;
    mem['h0E00] <= 32'h00E787B3;
    mem['h0E01] <= 32'h00379793;
    mem['h0E02] <= 32'h00078713;
    mem['h0E03] <= 32'hFEE44783;
    mem['h0E04] <= 32'h00F707B3;
    mem['h0E05] <= 32'h07C00713;
    mem['h0E06] <= 32'h00F707B3;
    mem['h0E07] <= 32'h00078023;
    mem['h0E08] <= 32'h5B80006F;
    mem['h0E09] <= 32'hFEF44703;
    mem['h0E0A] <= 32'h00070793;
    mem['h0E0B] <= 32'h00279793;
    mem['h0E0C] <= 32'h00E787B3;
    mem['h0E0D] <= 32'h00379793;
    mem['h0E0E] <= 32'h00078713;
    mem['h0E0F] <= 32'hFEE44783;
    mem['h0E10] <= 32'h00F707B3;
    mem['h0E11] <= 32'h07C00713;
    mem['h0E12] <= 32'h00F707B3;
    mem['h0E13] <= 32'h00900713;
    mem['h0E14] <= 32'h00E78023;
    mem['h0E15] <= 32'h5840006F;
    mem['h0E16] <= 32'hFEF44783;
    mem['h0E17] <= 32'hFD442703;
    mem['h0E18] <= 32'h06F70063;
    mem['h0E19] <= 32'hFEF44703;
    mem['h0E1A] <= 32'hFD442783;
    mem['h0E1B] <= 32'h00278793;
    mem['h0E1C] <= 32'h04F70863;
    mem['h0E1D] <= 32'hFEF44703;
    mem['h0E1E] <= 32'hFD442783;
    mem['h0E1F] <= 32'h00478793;
    mem['h0E20] <= 32'h04F70063;
    mem['h0E21] <= 32'hFEF44703;
    mem['h0E22] <= 32'hFD442783;
    mem['h0E23] <= 32'h00178793;
    mem['h0E24] <= 32'h00F71A63;
    mem['h0E25] <= 32'hFEE44703;
    mem['h0E26] <= 32'hFD842783;
    mem['h0E27] <= 32'h00278793;
    mem['h0E28] <= 32'h02F70063;
    mem['h0E29] <= 32'hFEF44703;
    mem['h0E2A] <= 32'hFD442783;
    mem['h0E2B] <= 32'h00378793;
    mem['h0E2C] <= 32'h04F71063;
    mem['h0E2D] <= 32'hFEE44783;
    mem['h0E2E] <= 32'hFD842703;
    mem['h0E2F] <= 32'h02F71A63;
    mem['h0E30] <= 32'hFEF44703;
    mem['h0E31] <= 32'h00070793;
    mem['h0E32] <= 32'h00279793;
    mem['h0E33] <= 32'h00E787B3;
    mem['h0E34] <= 32'h00379793;
    mem['h0E35] <= 32'h00078713;
    mem['h0E36] <= 32'hFEE44783;
    mem['h0E37] <= 32'h00F707B3;
    mem['h0E38] <= 32'h07C00713;
    mem['h0E39] <= 32'h00F707B3;
    mem['h0E3A] <= 32'h00078023;
    mem['h0E3B] <= 32'h4EC0006F;
    mem['h0E3C] <= 32'hFEF44703;
    mem['h0E3D] <= 32'h00070793;
    mem['h0E3E] <= 32'h00279793;
    mem['h0E3F] <= 32'h00E787B3;
    mem['h0E40] <= 32'h00379793;
    mem['h0E41] <= 32'h00078713;
    mem['h0E42] <= 32'hFEE44783;
    mem['h0E43] <= 32'h00F707B3;
    mem['h0E44] <= 32'h07C00713;
    mem['h0E45] <= 32'h00F707B3;
    mem['h0E46] <= 32'h00900713;
    mem['h0E47] <= 32'h00E78023;
    mem['h0E48] <= 32'h4B80006F;
    mem['h0E49] <= 32'hFEE44703;
    mem['h0E4A] <= 32'hFD842783;
    mem['h0E4B] <= 32'h00278793;
    mem['h0E4C] <= 32'h02F70863;
    mem['h0E4D] <= 32'hFEF44783;
    mem['h0E4E] <= 32'hFD442703;
    mem['h0E4F] <= 32'h02F70263;
    mem['h0E50] <= 32'hFEF44703;
    mem['h0E51] <= 32'hFD442783;
    mem['h0E52] <= 32'h00278793;
    mem['h0E53] <= 32'h00F70A63;
    mem['h0E54] <= 32'hFEF44703;
    mem['h0E55] <= 32'hFD442783;
    mem['h0E56] <= 32'h00478793;
    mem['h0E57] <= 32'h02F71A63;
    mem['h0E58] <= 32'hFEF44703;
    mem['h0E59] <= 32'h00070793;
    mem['h0E5A] <= 32'h00279793;
    mem['h0E5B] <= 32'h00E787B3;
    mem['h0E5C] <= 32'h00379793;
    mem['h0E5D] <= 32'h00078713;
    mem['h0E5E] <= 32'hFEE44783;
    mem['h0E5F] <= 32'h00F707B3;
    mem['h0E60] <= 32'h07C00713;
    mem['h0E61] <= 32'h00F707B3;
    mem['h0E62] <= 32'h00078023;
    mem['h0E63] <= 32'h44C0006F;
    mem['h0E64] <= 32'hFEF44703;
    mem['h0E65] <= 32'h00070793;
    mem['h0E66] <= 32'h00279793;
    mem['h0E67] <= 32'h00E787B3;
    mem['h0E68] <= 32'h00379793;
    mem['h0E69] <= 32'h00078713;
    mem['h0E6A] <= 32'hFEE44783;
    mem['h0E6B] <= 32'h00F707B3;
    mem['h0E6C] <= 32'h07C00713;
    mem['h0E6D] <= 32'h00F707B3;
    mem['h0E6E] <= 32'h00900713;
    mem['h0E6F] <= 32'h00E78023;
    mem['h0E70] <= 32'h4180006F;
    mem['h0E71] <= 32'hFEE44703;
    mem['h0E72] <= 32'hFD842783;
    mem['h0E73] <= 32'h00278793;
    mem['h0E74] <= 32'h02F70863;
    mem['h0E75] <= 32'hFEF44703;
    mem['h0E76] <= 32'hFD442783;
    mem['h0E77] <= 32'h00278793;
    mem['h0E78] <= 32'h02F70063;
    mem['h0E79] <= 32'hFEF44703;
    mem['h0E7A] <= 32'hFD442783;
    mem['h0E7B] <= 32'h00278793;
    mem['h0E7C] <= 32'h04E7C063;
    mem['h0E7D] <= 32'hFEE44783;
    mem['h0E7E] <= 32'hFD842703;
    mem['h0E7F] <= 32'h02F71A63;
    mem['h0E80] <= 32'hFEF44703;
    mem['h0E81] <= 32'h00070793;
    mem['h0E82] <= 32'h00279793;
    mem['h0E83] <= 32'h00E787B3;
    mem['h0E84] <= 32'h00379793;
    mem['h0E85] <= 32'h00078713;
    mem['h0E86] <= 32'hFEE44783;
    mem['h0E87] <= 32'h00F707B3;
    mem['h0E88] <= 32'h07C00713;
    mem['h0E89] <= 32'h00F707B3;
    mem['h0E8A] <= 32'h00078023;
    mem['h0E8B] <= 32'h3AC0006F;
    mem['h0E8C] <= 32'hFEF44703;
    mem['h0E8D] <= 32'h00070793;
    mem['h0E8E] <= 32'h00279793;
    mem['h0E8F] <= 32'h00E787B3;
    mem['h0E90] <= 32'h00379793;
    mem['h0E91] <= 32'h00078713;
    mem['h0E92] <= 32'hFEE44783;
    mem['h0E93] <= 32'h00F707B3;
    mem['h0E94] <= 32'h07C00713;
    mem['h0E95] <= 32'h00F707B3;
    mem['h0E96] <= 32'h00900713;
    mem['h0E97] <= 32'h00E78023;
    mem['h0E98] <= 32'h3780006F;
    mem['h0E99] <= 32'hFEF44783;
    mem['h0E9A] <= 32'hFD442703;
    mem['h0E9B] <= 32'h06F70063;
    mem['h0E9C] <= 32'hFEF44703;
    mem['h0E9D] <= 32'hFD442783;
    mem['h0E9E] <= 32'h00278793;
    mem['h0E9F] <= 32'h04F70863;
    mem['h0EA0] <= 32'hFEF44703;
    mem['h0EA1] <= 32'hFD442783;
    mem['h0EA2] <= 32'h00478793;
    mem['h0EA3] <= 32'h04F70063;
    mem['h0EA4] <= 32'hFEF44703;
    mem['h0EA5] <= 32'hFD442783;
    mem['h0EA6] <= 32'h00178793;
    mem['h0EA7] <= 32'h00F71863;
    mem['h0EA8] <= 32'hFEE44783;
    mem['h0EA9] <= 32'hFD842703;
    mem['h0EAA] <= 32'h02F70263;
    mem['h0EAB] <= 32'hFEF44703;
    mem['h0EAC] <= 32'hFD442783;
    mem['h0EAD] <= 32'h00378793;
    mem['h0EAE] <= 32'h04F71263;
    mem['h0EAF] <= 32'hFEE44703;
    mem['h0EB0] <= 32'hFD842783;
    mem['h0EB1] <= 32'h00278793;
    mem['h0EB2] <= 32'h02F71A63;
    mem['h0EB3] <= 32'hFEF44703;
    mem['h0EB4] <= 32'h00070793;
    mem['h0EB5] <= 32'h00279793;
    mem['h0EB6] <= 32'h00E787B3;
    mem['h0EB7] <= 32'h00379793;
    mem['h0EB8] <= 32'h00078713;
    mem['h0EB9] <= 32'hFEE44783;
    mem['h0EBA] <= 32'h00F707B3;
    mem['h0EBB] <= 32'h07C00713;
    mem['h0EBC] <= 32'h00F707B3;
    mem['h0EBD] <= 32'h00078023;
    mem['h0EBE] <= 32'h2E00006F;
    mem['h0EBF] <= 32'hFEF44703;
    mem['h0EC0] <= 32'h00070793;
    mem['h0EC1] <= 32'h00279793;
    mem['h0EC2] <= 32'h00E787B3;
    mem['h0EC3] <= 32'h00379793;
    mem['h0EC4] <= 32'h00078713;
    mem['h0EC5] <= 32'hFEE44783;
    mem['h0EC6] <= 32'h00F707B3;
    mem['h0EC7] <= 32'h07C00713;
    mem['h0EC8] <= 32'h00F707B3;
    mem['h0EC9] <= 32'h00900713;
    mem['h0ECA] <= 32'h00E78023;
    mem['h0ECB] <= 32'h2AC0006F;
    mem['h0ECC] <= 32'hFEE44783;
    mem['h0ECD] <= 32'hFD842703;
    mem['h0ECE] <= 32'h04F70863;
    mem['h0ECF] <= 32'hFEF44783;
    mem['h0ED0] <= 32'hFD442703;
    mem['h0ED1] <= 32'h04F70263;
    mem['h0ED2] <= 32'hFEF44703;
    mem['h0ED3] <= 32'hFD442783;
    mem['h0ED4] <= 32'h00278793;
    mem['h0ED5] <= 32'h02F70A63;
    mem['h0ED6] <= 32'hFEF44703;
    mem['h0ED7] <= 32'hFD442783;
    mem['h0ED8] <= 32'h00478793;
    mem['h0ED9] <= 32'h02F70263;
    mem['h0EDA] <= 32'hFEF44703;
    mem['h0EDB] <= 32'hFD442783;
    mem['h0EDC] <= 32'h00378793;
    mem['h0EDD] <= 32'h04F71263;
    mem['h0EDE] <= 32'hFEE44703;
    mem['h0EDF] <= 32'hFD842783;
    mem['h0EE0] <= 32'h00278793;
    mem['h0EE1] <= 32'h02F71A63;
    mem['h0EE2] <= 32'hFEF44703;
    mem['h0EE3] <= 32'h00070793;
    mem['h0EE4] <= 32'h00279793;
    mem['h0EE5] <= 32'h00E787B3;
    mem['h0EE6] <= 32'h00379793;
    mem['h0EE7] <= 32'h00078713;
    mem['h0EE8] <= 32'hFEE44783;
    mem['h0EE9] <= 32'h00F707B3;
    mem['h0EEA] <= 32'h07C00713;
    mem['h0EEB] <= 32'h00F707B3;
    mem['h0EEC] <= 32'h00078023;
    mem['h0EED] <= 32'h2240006F;
    mem['h0EEE] <= 32'hFEF44703;
    mem['h0EEF] <= 32'h00070793;
    mem['h0EF0] <= 32'h00279793;
    mem['h0EF1] <= 32'h00E787B3;
    mem['h0EF2] <= 32'h00379793;
    mem['h0EF3] <= 32'h00078713;
    mem['h0EF4] <= 32'hFEE44783;
    mem['h0EF5] <= 32'h00F707B3;
    mem['h0EF6] <= 32'h07C00713;
    mem['h0EF7] <= 32'h00F707B3;
    mem['h0EF8] <= 32'h00900713;
    mem['h0EF9] <= 32'h00E78023;
    mem['h0EFA] <= 32'h1F00006F;
    mem['h0EFB] <= 32'hFEE44703;
    mem['h0EFC] <= 32'hFD842783;
    mem['h0EFD] <= 32'h00278793;
    mem['h0EFE] <= 32'h00F70863;
    mem['h0EFF] <= 32'hFEF44783;
    mem['h0F00] <= 32'hFD442703;
    mem['h0F01] <= 32'h02F71A63;
    mem['h0F02] <= 32'hFEF44703;
    mem['h0F03] <= 32'h00070793;
    mem['h0F04] <= 32'h00279793;
    mem['h0F05] <= 32'h00E787B3;
    mem['h0F06] <= 32'h00379793;
    mem['h0F07] <= 32'h00078713;
    mem['h0F08] <= 32'hFEE44783;
    mem['h0F09] <= 32'h00F707B3;
    mem['h0F0A] <= 32'h07C00713;
    mem['h0F0B] <= 32'h00F707B3;
    mem['h0F0C] <= 32'h00078023;
    mem['h0F0D] <= 32'h1A40006F;
    mem['h0F0E] <= 32'hFEF44703;
    mem['h0F0F] <= 32'h00070793;
    mem['h0F10] <= 32'h00279793;
    mem['h0F11] <= 32'h00E787B3;
    mem['h0F12] <= 32'h00379793;
    mem['h0F13] <= 32'h00078713;
    mem['h0F14] <= 32'hFEE44783;
    mem['h0F15] <= 32'h00F707B3;
    mem['h0F16] <= 32'h07C00713;
    mem['h0F17] <= 32'h00F707B3;
    mem['h0F18] <= 32'h00900713;
    mem['h0F19] <= 32'h00E78023;
    mem['h0F1A] <= 32'h1700006F;
    mem['h0F1B] <= 32'hFEE44783;
    mem['h0F1C] <= 32'hFD842703;
    mem['h0F1D] <= 32'h04F70063;
    mem['h0F1E] <= 32'hFEE44703;
    mem['h0F1F] <= 32'hFD842783;
    mem['h0F20] <= 32'h00278793;
    mem['h0F21] <= 32'h02F70863;
    mem['h0F22] <= 32'hFEF44783;
    mem['h0F23] <= 32'hFD442703;
    mem['h0F24] <= 32'h02F70263;
    mem['h0F25] <= 32'hFEF44703;
    mem['h0F26] <= 32'hFD442783;
    mem['h0F27] <= 32'h00278793;
    mem['h0F28] <= 32'h00F70A63;
    mem['h0F29] <= 32'hFEF44703;
    mem['h0F2A] <= 32'hFD442783;
    mem['h0F2B] <= 32'h00478793;
    mem['h0F2C] <= 32'h02F71A63;
    mem['h0F2D] <= 32'hFEF44703;
    mem['h0F2E] <= 32'h00070793;
    mem['h0F2F] <= 32'h00279793;
    mem['h0F30] <= 32'h00E787B3;
    mem['h0F31] <= 32'h00379793;
    mem['h0F32] <= 32'h00078713;
    mem['h0F33] <= 32'hFEE44783;
    mem['h0F34] <= 32'h00F707B3;
    mem['h0F35] <= 32'h07C00713;
    mem['h0F36] <= 32'h00F707B3;
    mem['h0F37] <= 32'h00078023;
    mem['h0F38] <= 32'h0F80006F;
    mem['h0F39] <= 32'hFEF44703;
    mem['h0F3A] <= 32'h00070793;
    mem['h0F3B] <= 32'h00279793;
    mem['h0F3C] <= 32'h00E787B3;
    mem['h0F3D] <= 32'h00379793;
    mem['h0F3E] <= 32'h00078713;
    mem['h0F3F] <= 32'hFEE44783;
    mem['h0F40] <= 32'h00F707B3;
    mem['h0F41] <= 32'h07C00713;
    mem['h0F42] <= 32'h00F707B3;
    mem['h0F43] <= 32'h00900713;
    mem['h0F44] <= 32'h00E78023;
    mem['h0F45] <= 32'h0C40006F;
    mem['h0F46] <= 32'hFEE44703;
    mem['h0F47] <= 32'hFD842783;
    mem['h0F48] <= 32'h00278793;
    mem['h0F49] <= 32'h04F70663;
    mem['h0F4A] <= 32'hFEF44783;
    mem['h0F4B] <= 32'hFD442703;
    mem['h0F4C] <= 32'h04F70063;
    mem['h0F4D] <= 32'hFEF44703;
    mem['h0F4E] <= 32'hFD442783;
    mem['h0F4F] <= 32'h00278793;
    mem['h0F50] <= 32'h02F70863;
    mem['h0F51] <= 32'hFEF44703;
    mem['h0F52] <= 32'hFD442783;
    mem['h0F53] <= 32'h00478793;
    mem['h0F54] <= 32'h02F70063;
    mem['h0F55] <= 32'hFEF44703;
    mem['h0F56] <= 32'hFD442783;
    mem['h0F57] <= 32'h00178793;
    mem['h0F58] <= 32'h04F71063;
    mem['h0F59] <= 32'hFEE44783;
    mem['h0F5A] <= 32'hFD842703;
    mem['h0F5B] <= 32'h02F71A63;
    mem['h0F5C] <= 32'hFEF44703;
    mem['h0F5D] <= 32'h00070793;
    mem['h0F5E] <= 32'h00279793;
    mem['h0F5F] <= 32'h00E787B3;
    mem['h0F60] <= 32'h00379793;
    mem['h0F61] <= 32'h00078713;
    mem['h0F62] <= 32'hFEE44783;
    mem['h0F63] <= 32'h00F707B3;
    mem['h0F64] <= 32'h07C00713;
    mem['h0F65] <= 32'h00F707B3;
    mem['h0F66] <= 32'h00078023;
    mem['h0F67] <= 32'h03C0006F;
    mem['h0F68] <= 32'hFEF44703;
    mem['h0F69] <= 32'h00070793;
    mem['h0F6A] <= 32'h00279793;
    mem['h0F6B] <= 32'h00E787B3;
    mem['h0F6C] <= 32'h00379793;
    mem['h0F6D] <= 32'h00078713;
    mem['h0F6E] <= 32'hFEE44783;
    mem['h0F6F] <= 32'h00F707B3;
    mem['h0F70] <= 32'h07C00713;
    mem['h0F71] <= 32'h00F707B3;
    mem['h0F72] <= 32'h00900713;
    mem['h0F73] <= 32'h00E78023;
    mem['h0F74] <= 32'h0080006F;
    mem['h0F75] <= 32'h00000013;
    mem['h0F76] <= 32'hFEE44783;
    mem['h0F77] <= 32'h00178793;
    mem['h0F78] <= 32'hFEF40723;
    mem['h0F79] <= 32'hFD842783;
    mem['h0F7A] <= 32'h00278713;
    mem['h0F7B] <= 32'hFEE44783;
    mem['h0F7C] <= 32'h92F750E3;
    mem['h0F7D] <= 32'hFEF44783;
    mem['h0F7E] <= 32'h00178793;
    mem['h0F7F] <= 32'hFEF407A3;
    mem['h0F80] <= 32'hFD442783;
    mem['h0F81] <= 32'h00478713;
    mem['h0F82] <= 32'hFEF44783;
    mem['h0F83] <= 32'h8EF75CE3;
    mem['h0F84] <= 32'h00000013;
    mem['h0F85] <= 32'h00000013;
    mem['h0F86] <= 32'h02C12403;
    mem['h0F87] <= 32'h03010113;
    mem['h0F88] <= 32'h00008067;
    mem['h0F89] <= 32'hFC010113;
    mem['h0F8A] <= 32'h02112E23;
    mem['h0F8B] <= 32'h02812C23;
    mem['h0F8C] <= 32'h04010413;
    mem['h0F8D] <= 32'hFCA42623;
    mem['h0F8E] <= 32'hFCB42423;
    mem['h0F8F] <= 32'hFCC42223;
    mem['h0F90] <= 32'hFC042E23;
    mem['h0F91] <= 32'hFE042023;
    mem['h0F92] <= 32'hFE042223;
    mem['h0F93] <= 32'hFE042423;
    mem['h0F94] <= 32'hFE042623;
    mem['h0F95] <= 32'h03C0006F;
    mem['h0F96] <= 32'hFEC42783;
    mem['h0F97] <= 32'h00178713;
    mem['h0F98] <= 32'hFEE42623;
    mem['h0F99] <= 32'hFCC42683;
    mem['h0F9A] <= 32'h00A00713;
    mem['h0F9B] <= 32'h02E6E733;
    mem['h0F9C] <= 32'h00279793;
    mem['h0F9D] <= 32'hFF040693;
    mem['h0F9E] <= 32'h00F687B3;
    mem['h0F9F] <= 32'hFEE7A623;
    mem['h0FA0] <= 32'hFCC42703;
    mem['h0FA1] <= 32'h00A00793;
    mem['h0FA2] <= 32'h02F747B3;
    mem['h0FA3] <= 32'hFCF42623;
    mem['h0FA4] <= 32'hFCC42783;
    mem['h0FA5] <= 32'hFC0792E3;
    mem['h0FA6] <= 32'h00300793;
    mem['h0FA7] <= 32'hFEF42623;
    mem['h0FA8] <= 32'h04C0006F;
    mem['h0FA9] <= 32'hFEC42783;
    mem['h0FAA] <= 32'h00279793;
    mem['h0FAB] <= 32'hFF040713;
    mem['h0FAC] <= 32'h00F707B3;
    mem['h0FAD] <= 32'hFEC7A683;
    mem['h0FAE] <= 32'h00300713;
    mem['h0FAF] <= 32'hFEC42783;
    mem['h0FB0] <= 32'h40F707B3;
    mem['h0FB1] <= 32'h00279713;
    mem['h0FB2] <= 32'hFC842783;
    mem['h0FB3] <= 32'h00F707B3;
    mem['h0FB4] <= 32'hFC442603;
    mem['h0FB5] <= 32'h00078593;
    mem['h0FB6] <= 32'h00068513;
    mem['h0FB7] <= 32'h805FF0EF;
    mem['h0FB8] <= 32'hFEC42783;
    mem['h0FB9] <= 32'hFFF78793;
    mem['h0FBA] <= 32'hFEF42623;
    mem['h0FBB] <= 32'hFEC42783;
    mem['h0FBC] <= 32'hFA07DAE3;
    mem['h0FBD] <= 32'h00000013;
    mem['h0FBE] <= 32'h00000013;
    mem['h0FBF] <= 32'h03C12083;
    mem['h0FC0] <= 32'h03812403;
    mem['h0FC1] <= 32'h04010113;
    mem['h0FC2] <= 32'h00008067;
    mem['h0FC3] <= 32'hFD010113;
    mem['h0FC4] <= 32'h02112623;
    mem['h0FC5] <= 32'h02812423;
    mem['h0FC6] <= 32'h03010413;
    mem['h0FC7] <= 32'hFCA42E23;
    mem['h0FC8] <= 32'h01800793;
    mem['h0FC9] <= 32'hFEF407A3;
    mem['h0FCA] <= 32'h4600006F;
    mem['h0FCB] <= 32'h00300793;
    mem['h0FCC] <= 32'hFEF40723;
    mem['h0FCD] <= 32'h43C0006F;
    mem['h0FCE] <= 32'hFEE44703;
    mem['h0FCF] <= 32'h00300793;
    mem['h0FD0] <= 32'h00F70863;
    mem['h0FD1] <= 32'hFEE44703;
    mem['h0FD2] <= 32'h00400793;
    mem['h0FD3] <= 32'h0AF71E63;
    mem['h0FD4] <= 32'hFEF44703;
    mem['h0FD5] <= 32'h01800793;
    mem['h0FD6] <= 32'h04F70663;
    mem['h0FD7] <= 32'hFEF44703;
    mem['h0FD8] <= 32'h01A00793;
    mem['h0FD9] <= 32'h04F70063;
    mem['h0FDA] <= 32'hFEF44703;
    mem['h0FDB] <= 32'h01C00793;
    mem['h0FDC] <= 32'h02F70A63;
    mem['h0FDD] <= 32'hFEE44703;
    mem['h0FDE] <= 32'h00300793;
    mem['h0FDF] <= 32'h00F71863;
    mem['h0FE0] <= 32'hFEF44703;
    mem['h0FE1] <= 32'h01900793;
    mem['h0FE2] <= 32'h00F70E63;
    mem['h0FE3] <= 32'hFEE44703;
    mem['h0FE4] <= 32'h00400793;
    mem['h0FE5] <= 32'h04F71063;
    mem['h0FE6] <= 32'hFEF44703;
    mem['h0FE7] <= 32'h01B00793;
    mem['h0FE8] <= 32'h02F71A63;
    mem['h0FE9] <= 32'hFEF44703;
    mem['h0FEA] <= 32'h00070793;
    mem['h0FEB] <= 32'h00279793;
    mem['h0FEC] <= 32'h00E787B3;
    mem['h0FED] <= 32'h00379793;
    mem['h0FEE] <= 32'h00078713;
    mem['h0FEF] <= 32'hFEE44783;
    mem['h0FF0] <= 32'h00F707B3;
    mem['h0FF1] <= 32'h07C00713;
    mem['h0FF2] <= 32'h00F707B3;
    mem['h0FF3] <= 32'h00078023;
    mem['h0FF4] <= 32'h3940006F;
    mem['h0FF5] <= 32'hFEF44703;
    mem['h0FF6] <= 32'h00070793;
    mem['h0FF7] <= 32'h00279793;
    mem['h0FF8] <= 32'h00E787B3;
    mem['h0FF9] <= 32'h00379793;
    mem['h0FFA] <= 32'h00078713;
    mem['h0FFB] <= 32'hFEE44783;
    mem['h0FFC] <= 32'h00F707B3;
    mem['h0FFD] <= 32'h07C00713;
    mem['h0FFE] <= 32'h00F707B3;
    mem['h0FFF] <= 32'h00900713;
    mem['h1000] <= 32'h00E78023;
    mem['h1001] <= 32'h3600006F;
    mem['h1002] <= 32'hFEE44703;
    mem['h1003] <= 32'h00600793;
    mem['h1004] <= 32'h00F70863;
    mem['h1005] <= 32'hFEE44703;
    mem['h1006] <= 32'h00700793;
    mem['h1007] <= 32'h08F71663;
    mem['h1008] <= 32'hFEE44703;
    mem['h1009] <= 32'h00600793;
    mem['h100A] <= 32'h00F70E63;
    mem['h100B] <= 32'hFEF44703;
    mem['h100C] <= 32'h01800793;
    mem['h100D] <= 32'h00F70863;
    mem['h100E] <= 32'hFEF44703;
    mem['h100F] <= 32'h01C00793;
    mem['h1010] <= 32'h02F71A63;
    mem['h1011] <= 32'hFEF44703;
    mem['h1012] <= 32'h00070793;
    mem['h1013] <= 32'h00279793;
    mem['h1014] <= 32'h00E787B3;
    mem['h1015] <= 32'h00379793;
    mem['h1016] <= 32'h00078713;
    mem['h1017] <= 32'hFEE44783;
    mem['h1018] <= 32'h00F707B3;
    mem['h1019] <= 32'h07C00713;
    mem['h101A] <= 32'h00F707B3;
    mem['h101B] <= 32'h00078023;
    mem['h101C] <= 32'h2F40006F;
    mem['h101D] <= 32'hFEF44703;
    mem['h101E] <= 32'h00070793;
    mem['h101F] <= 32'h00279793;
    mem['h1020] <= 32'h00E787B3;
    mem['h1021] <= 32'h00379793;
    mem['h1022] <= 32'h00078713;
    mem['h1023] <= 32'hFEE44783;
    mem['h1024] <= 32'h00F707B3;
    mem['h1025] <= 32'h07C00713;
    mem['h1026] <= 32'h00F707B3;
    mem['h1027] <= 32'h00900713;
    mem['h1028] <= 32'h00E78023;
    mem['h1029] <= 32'h2C00006F;
    mem['h102A] <= 32'hFEE44703;
    mem['h102B] <= 32'h00900793;
    mem['h102C] <= 32'h00F70E63;
    mem['h102D] <= 32'hFEE44703;
    mem['h102E] <= 32'h00A00793;
    mem['h102F] <= 32'h00F70863;
    mem['h1030] <= 32'hFEE44703;
    mem['h1031] <= 32'h00B00793;
    mem['h1032] <= 32'h08F71C63;
    mem['h1033] <= 32'hFEE44703;
    mem['h1034] <= 32'h00900793;
    mem['h1035] <= 32'h02F70463;
    mem['h1036] <= 32'hFEE44703;
    mem['h1037] <= 32'h00B00793;
    mem['h1038] <= 32'h00F70E63;
    mem['h1039] <= 32'hFEF44703;
    mem['h103A] <= 32'h01800793;
    mem['h103B] <= 32'h00F70863;
    mem['h103C] <= 32'hFEF44703;
    mem['h103D] <= 32'h01C00793;
    mem['h103E] <= 32'h02F71A63;
    mem['h103F] <= 32'hFEF44703;
    mem['h1040] <= 32'h00070793;
    mem['h1041] <= 32'h00279793;
    mem['h1042] <= 32'h00E787B3;
    mem['h1043] <= 32'h00379793;
    mem['h1044] <= 32'h00078713;
    mem['h1045] <= 32'hFEE44783;
    mem['h1046] <= 32'h00F707B3;
    mem['h1047] <= 32'h07C00713;
    mem['h1048] <= 32'h00F707B3;
    mem['h1049] <= 32'h00078023;
    mem['h104A] <= 32'h23C0006F;
    mem['h104B] <= 32'hFEF44703;
    mem['h104C] <= 32'h00070793;
    mem['h104D] <= 32'h00279793;
    mem['h104E] <= 32'h00E787B3;
    mem['h104F] <= 32'h00379793;
    mem['h1050] <= 32'h00078713;
    mem['h1051] <= 32'hFEE44783;
    mem['h1052] <= 32'h00F707B3;
    mem['h1053] <= 32'h07C00713;
    mem['h1054] <= 32'h00F707B3;
    mem['h1055] <= 32'h00900713;
    mem['h1056] <= 32'h00E78023;
    mem['h1057] <= 32'h2080006F;
    mem['h1058] <= 32'hFEE44703;
    mem['h1059] <= 32'h00D00793;
    mem['h105A] <= 32'h00F70E63;
    mem['h105B] <= 32'hFEE44703;
    mem['h105C] <= 32'h00E00793;
    mem['h105D] <= 32'h00F70863;
    mem['h105E] <= 32'hFEE44703;
    mem['h105F] <= 32'h00F00793;
    mem['h1060] <= 32'h0AF71E63;
    mem['h1061] <= 32'hFEE44703;
    mem['h1062] <= 32'h00D00793;
    mem['h1063] <= 32'h04F70663;
    mem['h1064] <= 32'hFEE44703;
    mem['h1065] <= 32'h00E00793;
    mem['h1066] <= 32'h00F71E63;
    mem['h1067] <= 32'hFEF44703;
    mem['h1068] <= 32'h01800793;
    mem['h1069] <= 32'h02F70A63;
    mem['h106A] <= 32'hFEF44703;
    mem['h106B] <= 32'h01A00793;
    mem['h106C] <= 32'h02F70463;
    mem['h106D] <= 32'hFEE44703;
    mem['h106E] <= 32'h00F00793;
    mem['h106F] <= 32'h04F71663;
    mem['h1070] <= 32'hFEF44703;
    mem['h1071] <= 32'h01900793;
    mem['h1072] <= 32'h00F70863;
    mem['h1073] <= 32'hFEF44703;
    mem['h1074] <= 32'h01A00793;
    mem['h1075] <= 32'h02E7FA63;
    mem['h1076] <= 32'hFEF44703;
    mem['h1077] <= 32'h00070793;
    mem['h1078] <= 32'h00279793;
    mem['h1079] <= 32'h00E787B3;
    mem['h107A] <= 32'h00379793;
    mem['h107B] <= 32'h00078713;
    mem['h107C] <= 32'hFEE44783;
    mem['h107D] <= 32'h00F707B3;
    mem['h107E] <= 32'h07C00713;
    mem['h107F] <= 32'h00F707B3;
    mem['h1080] <= 32'h00078023;
    mem['h1081] <= 32'h1600006F;
    mem['h1082] <= 32'hFEF44703;
    mem['h1083] <= 32'h00070793;
    mem['h1084] <= 32'h00279793;
    mem['h1085] <= 32'h00E787B3;
    mem['h1086] <= 32'h00379793;
    mem['h1087] <= 32'h00078713;
    mem['h1088] <= 32'hFEE44783;
    mem['h1089] <= 32'h00F707B3;
    mem['h108A] <= 32'h07C00713;
    mem['h108B] <= 32'h00F707B3;
    mem['h108C] <= 32'h00900713;
    mem['h108D] <= 32'h00E78023;
    mem['h108E] <= 32'h12C0006F;
    mem['h108F] <= 32'hFEE44703;
    mem['h1090] <= 32'h01100793;
    mem['h1091] <= 32'h00F70863;
    mem['h1092] <= 32'hFEE44703;
    mem['h1093] <= 32'h01200793;
    mem['h1094] <= 32'h08F71863;
    mem['h1095] <= 32'hFEE44703;
    mem['h1096] <= 32'h01100793;
    mem['h1097] <= 32'h02F70063;
    mem['h1098] <= 32'hFEE44703;
    mem['h1099] <= 32'h01200793;
    mem['h109A] <= 32'h04F71263;
    mem['h109B] <= 32'hFEF44783;
    mem['h109C] <= 32'h0017F793;
    mem['h109D] <= 32'h0FF7F793;
    mem['h109E] <= 32'h02079A63;
    mem['h109F] <= 32'hFEF44703;
    mem['h10A0] <= 32'h00070793;
    mem['h10A1] <= 32'h00279793;
    mem['h10A2] <= 32'h00E787B3;
    mem['h10A3] <= 32'h00379793;
    mem['h10A4] <= 32'h00078713;
    mem['h10A5] <= 32'hFEE44783;
    mem['h10A6] <= 32'h00F707B3;
    mem['h10A7] <= 32'h07C00713;
    mem['h10A8] <= 32'h00F707B3;
    mem['h10A9] <= 32'h00078023;
    mem['h10AA] <= 32'h0BC0006F;
    mem['h10AB] <= 32'hFEF44703;
    mem['h10AC] <= 32'h00070793;
    mem['h10AD] <= 32'h00279793;
    mem['h10AE] <= 32'h00E787B3;
    mem['h10AF] <= 32'h00379793;
    mem['h10B0] <= 32'h00078713;
    mem['h10B1] <= 32'hFEE44783;
    mem['h10B2] <= 32'h00F707B3;
    mem['h10B3] <= 32'h07C00713;
    mem['h10B4] <= 32'h00F707B3;
    mem['h10B5] <= 32'h00900713;
    mem['h10B6] <= 32'h00E78023;
    mem['h10B7] <= 32'h0880006F;
    mem['h10B8] <= 32'hFEE44703;
    mem['h10B9] <= 32'h01400793;
    mem['h10BA] <= 32'h06F71E63;
    mem['h10BB] <= 32'hFEF44703;
    mem['h10BC] <= 32'h01900793;
    mem['h10BD] <= 32'h00F70863;
    mem['h10BE] <= 32'hFEF44703;
    mem['h10BF] <= 32'h01B00793;
    mem['h10C0] <= 32'h02F71A63;
    mem['h10C1] <= 32'hFEF44703;
    mem['h10C2] <= 32'h00070793;
    mem['h10C3] <= 32'h00279793;
    mem['h10C4] <= 32'h00E787B3;
    mem['h10C5] <= 32'h00379793;
    mem['h10C6] <= 32'h00078713;
    mem['h10C7] <= 32'hFEE44783;
    mem['h10C8] <= 32'h00F707B3;
    mem['h10C9] <= 32'h07C00713;
    mem['h10CA] <= 32'h00F707B3;
    mem['h10CB] <= 32'h00078023;
    mem['h10CC] <= 32'h0340006F;
    mem['h10CD] <= 32'hFEF44703;
    mem['h10CE] <= 32'h00070793;
    mem['h10CF] <= 32'h00279793;
    mem['h10D0] <= 32'h00E787B3;
    mem['h10D1] <= 32'h00379793;
    mem['h10D2] <= 32'h00078713;
    mem['h10D3] <= 32'hFEE44783;
    mem['h10D4] <= 32'h00F707B3;
    mem['h10D5] <= 32'h07C00713;
    mem['h10D6] <= 32'h00F707B3;
    mem['h10D7] <= 32'h00900713;
    mem['h10D8] <= 32'h00E78023;
    mem['h10D9] <= 32'hFEE44783;
    mem['h10DA] <= 32'h00178793;
    mem['h10DB] <= 32'hFEF40723;
    mem['h10DC] <= 32'hFEE44703;
    mem['h10DD] <= 32'h01400793;
    mem['h10DE] <= 32'hBCE7F0E3;
    mem['h10DF] <= 32'hFEF44783;
    mem['h10E0] <= 32'h00178793;
    mem['h10E1] <= 32'hFEF407A3;
    mem['h10E2] <= 32'hFEF44703;
    mem['h10E3] <= 32'h01C00793;
    mem['h10E4] <= 32'hB8E7FEE3;
    mem['h10E5] <= 32'h01800613;
    mem['h10E6] <= 32'h01600593;
    mem['h10E7] <= 32'hFDC42503;
    mem['h10E8] <= 32'hA85FF0EF;
    mem['h10E9] <= 32'h00000013;
    mem['h10EA] <= 32'h02C12083;
    mem['h10EB] <= 32'h02812403;
    mem['h10EC] <= 32'h03010113;
    mem['h10ED] <= 32'h00008067;
    mem['h10EE] <= 32'hFE010113;
    mem['h10EF] <= 32'h00812E23;
    mem['h10F0] <= 32'h02010413;
    mem['h10F1] <= 32'hFE0407A3;
    mem['h10F2] <= 32'h0940006F;
    mem['h10F3] <= 32'hFE040723;
    mem['h10F4] <= 32'h0740006F;
    mem['h10F5] <= 32'hFEF44783;
    mem['h10F6] <= 32'h02078463;
    mem['h10F7] <= 32'hFEF44703;
    mem['h10F8] <= 32'h01600793;
    mem['h10F9] <= 32'h00E7EE63;
    mem['h10FA] <= 32'hFEE44703;
    mem['h10FB] <= 32'h01300793;
    mem['h10FC] <= 32'h00F70863;
    mem['h10FD] <= 32'hFEE44703;
    mem['h10FE] <= 32'h01400793;
    mem['h10FF] <= 32'h00F71663;
    mem['h1100] <= 32'h00900713;
    mem['h1101] <= 32'h0080006F;
    mem['h1102] <= 32'h00000713;
    mem['h1103] <= 32'hFEF44683;
    mem['h1104] <= 32'h00068793;
    mem['h1105] <= 32'h00279793;
    mem['h1106] <= 32'h00D787B3;
    mem['h1107] <= 32'h00379793;
    mem['h1108] <= 32'h00078693;
    mem['h1109] <= 32'hFEE44783;
    mem['h110A] <= 32'h00F687B3;
    mem['h110B] <= 32'h07C00693;
    mem['h110C] <= 32'h00F687B3;
    mem['h110D] <= 32'h00E78023;
    mem['h110E] <= 32'hFEE44783;
    mem['h110F] <= 32'h00178793;
    mem['h1110] <= 32'hFEF40723;
    mem['h1111] <= 32'hFEE44703;
    mem['h1112] <= 32'h02700793;
    mem['h1113] <= 32'hF8E7F4E3;
    mem['h1114] <= 32'hFEF44783;
    mem['h1115] <= 32'h00178793;
    mem['h1116] <= 32'hFEF407A3;
    mem['h1117] <= 32'hFEF44703;
    mem['h1118] <= 32'h01D00793;
    mem['h1119] <= 32'hF6E7F4E3;
    mem['h111A] <= 32'h00000013;
    mem['h111B] <= 32'h00000013;
    mem['h111C] <= 32'h01C12403;
    mem['h111D] <= 32'h02010113;
    mem['h111E] <= 32'h00008067;
    mem['h111F] <= 32'hFD010113;
    mem['h1120] <= 32'h02112623;
    mem['h1121] <= 32'h02812423;
    mem['h1122] <= 32'h03010413;
    mem['h1123] <= 32'hFCA42E23;
    mem['h1124] <= 32'hFE041723;
    mem['h1125] <= 32'hFE042423;
    mem['h1126] <= 32'h0340006F;
    mem['h1127] <= 32'h001057B7;
    mem['h1128] <= 32'h48478513;
    mem['h1129] <= 32'h6E9000EF;
    mem['h112A] <= 32'hFE842783;
    mem['h112B] <= 32'h0017F793;
    mem['h112C] <= 32'h00079863;
    mem['h112D] <= 32'hFEE45783;
    mem['h112E] <= 32'h00178793;
    mem['h112F] <= 32'hFEF41723;
    mem['h1130] <= 32'hFE842783;
    mem['h1131] <= 32'h00178793;
    mem['h1132] <= 32'hFEF42423;
    mem['h1133] <= 32'hFE842703;
    mem['h1134] <= 32'hFDC42783;
    mem['h1135] <= 32'hFCF764E3;
    mem['h1136] <= 32'h00000013;
    mem['h1137] <= 32'h00000013;
    mem['h1138] <= 32'h02C12083;
    mem['h1139] <= 32'h02812403;
    mem['h113A] <= 32'h03010113;
    mem['h113B] <= 32'h00008067;
    mem['h113C] <= 32'hFD010113;
    mem['h113D] <= 32'h02812623;
    mem['h113E] <= 32'h03010413;
    mem['h113F] <= 32'hFCA42E23;
    mem['h1140] <= 32'hFDC42783;
    mem['h1141] <= 32'h0007A783;
    mem['h1142] <= 32'hFEF42623;
    mem['h1143] <= 32'hFEC42783;
    mem['h1144] <= 32'h00D79793;
    mem['h1145] <= 32'hFEC42703;
    mem['h1146] <= 32'h00F747B3;
    mem['h1147] <= 32'hFEF42623;
    mem['h1148] <= 32'hFEC42783;
    mem['h1149] <= 32'h0117D793;
    mem['h114A] <= 32'hFEC42703;
    mem['h114B] <= 32'h00F747B3;
    mem['h114C] <= 32'hFEF42623;
    mem['h114D] <= 32'hFEC42783;
    mem['h114E] <= 32'h00579793;
    mem['h114F] <= 32'hFEC42703;
    mem['h1150] <= 32'h00F747B3;
    mem['h1151] <= 32'hFEF42623;
    mem['h1152] <= 32'hFDC42783;
    mem['h1153] <= 32'hFEC42703;
    mem['h1154] <= 32'h00E7A023;
    mem['h1155] <= 32'hFEC42783;
    mem['h1156] <= 32'h00078513;
    mem['h1157] <= 32'h02C12403;
    mem['h1158] <= 32'h03010113;
    mem['h1159] <= 32'h00008067;
    mem['h115A] <= 32'hFF010113;
    mem['h115B] <= 32'h00112623;
    mem['h115C] <= 32'h00812423;
    mem['h115D] <= 32'h01010413;
    mem['h115E] <= 32'h07400513;
    mem['h115F] <= 32'hF75FF0EF;
    mem['h1160] <= 32'h00050793;
    mem['h1161] <= 32'h0017F793;
    mem['h1162] <= 32'h00078513;
    mem['h1163] <= 32'h00C12083;
    mem['h1164] <= 32'h00812403;
    mem['h1165] <= 32'h01010113;
    mem['h1166] <= 32'h00008067;
    mem['h1167] <= 32'hFD010113;
    mem['h1168] <= 32'h02112623;
    mem['h1169] <= 32'h02812423;
    mem['h116A] <= 32'h03010413;
    mem['h116B] <= 32'hFCA42E23;
    mem['h116C] <= 32'hFCB42C23;
    mem['h116D] <= 32'hFD842703;
    mem['h116E] <= 32'hFDC42783;
    mem['h116F] <= 32'h40F707B3;
    mem['h1170] <= 32'h00178793;
    mem['h1171] <= 32'hFEF42623;
    mem['h1172] <= 32'h07800513;
    mem['h1173] <= 32'hF25FF0EF;
    mem['h1174] <= 32'h00050713;
    mem['h1175] <= 32'hFEC42783;
    mem['h1176] <= 32'h02F77733;
    mem['h1177] <= 32'hFDC42783;
    mem['h1178] <= 32'h00F707B3;
    mem['h1179] <= 32'hFEF42423;
    mem['h117A] <= 32'hFE842783;
    mem['h117B] <= 32'h00078513;
    mem['h117C] <= 32'h02C12083;
    mem['h117D] <= 32'h02812403;
    mem['h117E] <= 32'h03010113;
    mem['h117F] <= 32'h00008067;
    mem['h1180] <= 32'hF9010113;
    mem['h1181] <= 32'h06112623;
    mem['h1182] <= 32'h06812423;
    mem['h1183] <= 32'h06912223;
    mem['h1184] <= 32'h07010413;
    mem['h1185] <= 32'h020007B7;
    mem['h1186] <= 32'h00478793;
    mem['h1187] <= 32'h0D900713;
    mem['h1188] <= 32'h00E7A023;
    mem['h1189] <= 32'h001057B7;
    mem['h118A] <= 32'h49478513;
    mem['h118B] <= 32'h561000EF;
    mem['h118C] <= 32'hFE0407A3;
    mem['h118D] <= 32'hFE040723;
    mem['h118E] <= 32'hFE0406A3;
    mem['h118F] <= 32'hFE040623;
    mem['h1190] <= 32'hFE0405A3;
    mem['h1191] <= 32'h030007B7;
    mem['h1192] <= 32'h0007A023;
    mem['h1193] <= 32'h955FE0EF;
    mem['h1194] <= 32'hAB5FB0EF;
    mem['h1195] <= 32'h000017B7;
    mem['h1196] <= 32'hBB878513;
    mem['h1197] <= 32'hE21FF0EF;
    mem['h1198] <= 32'hF85FB0EF;
    mem['h1199] <= 32'h000017B7;
    mem['h119A] <= 32'hBB878513;
    mem['h119B] <= 32'hE11FF0EF;
    mem['h119C] <= 32'h9C5FC0EF;
    mem['h119D] <= 32'h000017B7;
    mem['h119E] <= 32'hBB878513;
    mem['h119F] <= 32'hE01FF0EF;
    mem['h11A0] <= 32'hD39FF0EF;
    mem['h11A1] <= 32'h00900513;
    mem['h11A2] <= 32'hB0DFD0EF;
    mem['h11A3] <= 32'h00300613;
    mem['h11A4] <= 32'h00900593;
    mem['h11A5] <= 32'h00500513;
    mem['h11A6] <= 32'hC18FD0EF;
    mem['h11A7] <= 32'h00300613;
    mem['h11A8] <= 32'h00900593;
    mem['h11A9] <= 32'h00F00513;
    mem['h11AA] <= 32'hC08FD0EF;
    mem['h11AB] <= 32'h00300613;
    mem['h11AC] <= 32'h00900593;
    mem['h11AD] <= 32'h01900513;
    mem['h11AE] <= 32'hBF8FD0EF;
    mem['h11AF] <= 32'h000017B7;
    mem['h11B0] <= 32'hFA078513;
    mem['h11B1] <= 32'hDB9FF0EF;
    mem['h11B2] <= 32'hFE041423;
    mem['h11B3] <= 32'h00300793;
    mem['h11B4] <= 32'hFEF403A3;
    mem['h11B5] <= 32'hFE040323;
    mem['h11B6] <= 32'h00F00793;
    mem['h11B7] <= 32'hFEF402A3;
    mem['h11B8] <= 32'h00F00793;
    mem['h11B9] <= 32'hFEF40223;
    mem['h11BA] <= 32'hFE0401A3;
    mem['h11BB] <= 32'h00300793;
    mem['h11BC] <= 32'hFEF40123;
    mem['h11BD] <= 32'hFA0400A3;
    mem['h11BE] <= 32'h00100793;
    mem['h11BF] <= 32'hFEF400A3;
    mem['h11C0] <= 32'hFC041F23;
    mem['h11C1] <= 32'hFC041E23;
    mem['h11C2] <= 32'hF8042E23;
    mem['h11C3] <= 32'hFC040DA3;
    mem['h11C4] <= 32'hFC040D23;
    mem['h11C5] <= 32'hFC040CA3;
    mem['h11C6] <= 32'hFC040C23;
    mem['h11C7] <= 32'hFC040BA3;
    mem['h11C8] <= 32'hFC040B23;
    mem['h11C9] <= 32'hFDC45783;
    mem['h11CA] <= 32'h00078513;
    mem['h11CB] <= 32'hFE0FF0EF;
    mem['h11CC] <= 32'hFDA44783;
    mem['h11CD] <= 32'h00078E63;
    mem['h11CE] <= 32'hFE244703;
    mem['h11CF] <= 32'h00100793;
    mem['h11D0] <= 32'h00F71863;
    mem['h11D1] <= 32'h00100793;
    mem['h11D2] <= 32'hFCF40CA3;
    mem['h11D3] <= 32'hFC040D23;
    mem['h11D4] <= 32'hFDA44783;
    mem['h11D5] <= 32'h0C078E63;
    mem['h11D6] <= 32'hFE244783;
    mem['h11D7] <= 32'hFFF78793;
    mem['h11D8] <= 32'hFEF40123;
    mem['h11D9] <= 32'hFE244783;
    mem['h11DA] <= 32'h00078513;
    mem['h11DB] <= 32'hAC1FD0EF;
    mem['h11DC] <= 32'h000017B7;
    mem['h11DD] <= 32'hFA078513;
    mem['h11DE] <= 32'hD05FF0EF;
    mem['h11DF] <= 32'hFC040AA3;
    mem['h11E0] <= 32'h0940006F;
    mem['h11E1] <= 32'hFC040A23;
    mem['h11E2] <= 32'h0740006F;
    mem['h11E3] <= 32'hFD544783;
    mem['h11E4] <= 32'h02078463;
    mem['h11E5] <= 32'hFD544703;
    mem['h11E6] <= 32'h01600793;
    mem['h11E7] <= 32'h00E7EE63;
    mem['h11E8] <= 32'hFD444703;
    mem['h11E9] <= 32'h01300793;
    mem['h11EA] <= 32'h00F70863;
    mem['h11EB] <= 32'hFD444703;
    mem['h11EC] <= 32'h01400793;
    mem['h11ED] <= 32'h00F71663;
    mem['h11EE] <= 32'h00900713;
    mem['h11EF] <= 32'h0080006F;
    mem['h11F0] <= 32'h00000713;
    mem['h11F1] <= 32'hFD544683;
    mem['h11F2] <= 32'h00068793;
    mem['h11F3] <= 32'h00279793;
    mem['h11F4] <= 32'h00D787B3;
    mem['h11F5] <= 32'h00379793;
    mem['h11F6] <= 32'h00078693;
    mem['h11F7] <= 32'hFD444783;
    mem['h11F8] <= 32'h00F687B3;
    mem['h11F9] <= 32'h07C00693;
    mem['h11FA] <= 32'h00F687B3;
    mem['h11FB] <= 32'h00E78023;
    mem['h11FC] <= 32'hFD444783;
    mem['h11FD] <= 32'h00178793;
    mem['h11FE] <= 32'hFCF40A23;
    mem['h11FF] <= 32'hFD444703;
    mem['h1200] <= 32'h02700793;
    mem['h1201] <= 32'hF8E7F4E3;
    mem['h1202] <= 32'hFD544783;
    mem['h1203] <= 32'h00178793;
    mem['h1204] <= 32'hFCF40AA3;
    mem['h1205] <= 32'hFD544703;
    mem['h1206] <= 32'h01D00793;
    mem['h1207] <= 32'hF6E7F4E3;
    mem['h1208] <= 32'hFC040D23;
    mem['h1209] <= 32'hFDC45783;
    mem['h120A] <= 32'h00078513;
    mem['h120B] <= 32'hEE0FF0EF;
    mem['h120C] <= 32'hFD944783;
    mem['h120D] <= 32'h0C078E63;
    mem['h120E] <= 32'hA80FE0EF;
    mem['h120F] <= 32'h0080006F;
    mem['h1210] <= 32'h895FB0EF;
    mem['h1211] <= 32'h52C04783;
    mem['h1212] <= 32'h0107F793;
    mem['h1213] <= 32'hFE078AE3;
    mem['h1214] <= 32'hFC0409A3;
    mem['h1215] <= 32'h0940006F;
    mem['h1216] <= 32'hFC040923;
    mem['h1217] <= 32'h0740006F;
    mem['h1218] <= 32'hFD344783;
    mem['h1219] <= 32'h02078463;
    mem['h121A] <= 32'hFD344703;
    mem['h121B] <= 32'h01600793;
    mem['h121C] <= 32'h00E7EE63;
    mem['h121D] <= 32'hFD244703;
    mem['h121E] <= 32'h01300793;
    mem['h121F] <= 32'h00F70863;
    mem['h1220] <= 32'hFD244703;
    mem['h1221] <= 32'h01400793;
    mem['h1222] <= 32'h00F71663;
    mem['h1223] <= 32'h00900713;
    mem['h1224] <= 32'h0080006F;
    mem['h1225] <= 32'h00000713;
    mem['h1226] <= 32'hFD344683;
    mem['h1227] <= 32'h00068793;
    mem['h1228] <= 32'h00279793;
    mem['h1229] <= 32'h00D787B3;
    mem['h122A] <= 32'h00379793;
    mem['h122B] <= 32'h00078693;
    mem['h122C] <= 32'hFD244783;
    mem['h122D] <= 32'h00F687B3;
    mem['h122E] <= 32'h07C00693;
    mem['h122F] <= 32'h00F687B3;
    mem['h1230] <= 32'h00E78023;
    mem['h1231] <= 32'hFD244783;
    mem['h1232] <= 32'h00178793;
    mem['h1233] <= 32'hFCF40923;
    mem['h1234] <= 32'hFD244703;
    mem['h1235] <= 32'h02700793;
    mem['h1236] <= 32'hF8E7F4E3;
    mem['h1237] <= 32'hFD344783;
    mem['h1238] <= 32'h00178793;
    mem['h1239] <= 32'hFCF409A3;
    mem['h123A] <= 32'hFD344703;
    mem['h123B] <= 32'h01D00793;
    mem['h123C] <= 32'hF6E7F4E3;
    mem['h123D] <= 32'hFC040CA3;
    mem['h123E] <= 32'hFC041E23;
    mem['h123F] <= 32'h00F00793;
    mem['h1240] <= 32'hFEF40223;
    mem['h1241] <= 32'hFDC45783;
    mem['h1242] <= 32'h00078513;
    mem['h1243] <= 32'hE00FF0EF;
    mem['h1244] <= 32'h07002783;
    mem['h1245] <= 32'hFFF78713;
    mem['h1246] <= 32'h06E02823;
    mem['h1247] <= 32'hFB8FB0EF;
    mem['h1248] <= 32'h52C04783;
    mem['h1249] <= 32'h0017F793;
    mem['h124A] <= 32'h00078C63;
    mem['h124B] <= 32'h00100793;
    mem['h124C] <= 32'hFEF40623;
    mem['h124D] <= 32'h001057B7;
    mem['h124E] <= 32'h4A478513;
    mem['h124F] <= 32'h251000EF;
    mem['h1250] <= 32'h52C04783;
    mem['h1251] <= 32'h0087F793;
    mem['h1252] <= 32'h00078C63;
    mem['h1253] <= 32'h00100793;
    mem['h1254] <= 32'hFEF40723;
    mem['h1255] <= 32'h001057B7;
    mem['h1256] <= 32'h4B078513;
    mem['h1257] <= 32'h231000EF;
    mem['h1258] <= 32'h52C04783;
    mem['h1259] <= 32'h0027F793;
    mem['h125A] <= 32'h00078C63;
    mem['h125B] <= 32'h00100793;
    mem['h125C] <= 32'hFEF407A3;
    mem['h125D] <= 32'h001057B7;
    mem['h125E] <= 32'h4C078513;
    mem['h125F] <= 32'h211000EF;
    mem['h1260] <= 32'h52C04783;
    mem['h1261] <= 32'h0047F793;
    mem['h1262] <= 32'h00078C63;
    mem['h1263] <= 32'h00100793;
    mem['h1264] <= 32'hFEF405A3;
    mem['h1265] <= 32'h001057B7;
    mem['h1266] <= 32'h4D078513;
    mem['h1267] <= 32'h1F1000EF;
    mem['h1268] <= 32'h52C04783;
    mem['h1269] <= 32'h0107F793;
    mem['h126A] <= 32'h00078C63;
    mem['h126B] <= 32'h00100793;
    mem['h126C] <= 32'hFEF406A3;
    mem['h126D] <= 32'h001057B7;
    mem['h126E] <= 32'h4E078513;
    mem['h126F] <= 32'h1D1000EF;
    mem['h1270] <= 32'h52C04783;
    mem['h1271] <= 32'h1007E713;
    mem['h1272] <= 32'h030007B7;
    mem['h1273] <= 32'h00E7A023;
    mem['h1274] <= 32'h07002783;
    mem['h1275] <= 32'hD4079EE3;
    mem['h1276] <= 32'h00001737;
    mem['h1277] <= 32'h9C470713;
    mem['h1278] <= 32'h06E02823;
    mem['h1279] <= 32'hFE344783;
    mem['h127A] <= 32'h00178793;
    mem['h127B] <= 32'hFEF401A3;
    mem['h127C] <= 32'hFE344703;
    mem['h127D] <= 32'hFE444783;
    mem['h127E] <= 32'h40F707B3;
    mem['h127F] <= 32'h0017B793;
    mem['h1280] <= 32'hFAF400A3;
    mem['h1281] <= 32'hFD644783;
    mem['h1282] <= 32'h0E079663;
    mem['h1283] <= 32'hFEE44783;
    mem['h1284] <= 32'h02078A63;
    mem['h1285] <= 32'hFE845703;
    mem['h1286] <= 32'hFE744583;
    mem['h1287] <= 32'hFE644603;
    mem['h1288] <= 32'hFE544783;
    mem['h1289] <= 32'h00178793;
    mem['h128A] <= 32'h00078693;
    mem['h128B] <= 32'h00070513;
    mem['h128C] <= 32'hB6DFE0EF;
    mem['h128D] <= 32'h00050793;
    mem['h128E] <= 32'h00078663;
    mem['h128F] <= 32'h00100793;
    mem['h1290] <= 32'h0080006F;
    mem['h1291] <= 32'h00000793;
    mem['h1292] <= 32'h0FF7F713;
    mem['h1293] <= 32'hFE544783;
    mem['h1294] <= 32'h00F707B3;
    mem['h1295] <= 32'hFEF402A3;
    mem['h1296] <= 32'hFEC44783;
    mem['h1297] <= 32'h02078A63;
    mem['h1298] <= 32'hFE845703;
    mem['h1299] <= 32'hFE744583;
    mem['h129A] <= 32'hFE644603;
    mem['h129B] <= 32'hFE544783;
    mem['h129C] <= 32'hFFF78793;
    mem['h129D] <= 32'h00078693;
    mem['h129E] <= 32'h00070513;
    mem['h129F] <= 32'hB21FE0EF;
    mem['h12A0] <= 32'h00050793;
    mem['h12A1] <= 32'h00078663;
    mem['h12A2] <= 32'h00100793;
    mem['h12A3] <= 32'h0080006F;
    mem['h12A4] <= 32'h00000793;
    mem['h12A5] <= 32'h0FF7F793;
    mem['h12A6] <= 32'hFE544703;
    mem['h12A7] <= 32'h40F707B3;
    mem['h12A8] <= 32'hFEF402A3;
    mem['h12A9] <= 32'hFEF44783;
    mem['h12AA] <= 32'h02078A63;
    mem['h12AB] <= 32'hFE845703;
    mem['h12AC] <= 32'hFE744583;
    mem['h12AD] <= 32'hFE644783;
    mem['h12AE] <= 32'h00178793;
    mem['h12AF] <= 32'hFE544683;
    mem['h12B0] <= 32'h00078613;
    mem['h12B1] <= 32'h00070513;
    mem['h12B2] <= 32'hAD5FE0EF;
    mem['h12B3] <= 32'h00050793;
    mem['h12B4] <= 32'h00078663;
    mem['h12B5] <= 32'h00100793;
    mem['h12B6] <= 32'h0080006F;
    mem['h12B7] <= 32'h00000793;
    mem['h12B8] <= 32'h0FF7F713;
    mem['h12B9] <= 32'hFE644783;
    mem['h12BA] <= 32'h00F707B3;
    mem['h12BB] <= 32'hFEF40323;
    mem['h12BC] <= 32'h0E80006F;
    mem['h12BD] <= 32'hFEC44783;
    mem['h12BE] <= 32'h02078A63;
    mem['h12BF] <= 32'hFE845703;
    mem['h12C0] <= 32'hFE744583;
    mem['h12C1] <= 32'hFE644603;
    mem['h12C2] <= 32'hFE544783;
    mem['h12C3] <= 32'hFFF78793;
    mem['h12C4] <= 32'h00078693;
    mem['h12C5] <= 32'h00070513;
    mem['h12C6] <= 32'hA85FE0EF;
    mem['h12C7] <= 32'h00050793;
    mem['h12C8] <= 32'h00078663;
    mem['h12C9] <= 32'h00100793;
    mem['h12CA] <= 32'h0080006F;
    mem['h12CB] <= 32'h00000793;
    mem['h12CC] <= 32'h0FF7F793;
    mem['h12CD] <= 32'hFE544703;
    mem['h12CE] <= 32'h40F707B3;
    mem['h12CF] <= 32'hFEF402A3;
    mem['h12D0] <= 32'hFEE44783;
    mem['h12D1] <= 32'h02078A63;
    mem['h12D2] <= 32'hFE845703;
    mem['h12D3] <= 32'hFE744583;
    mem['h12D4] <= 32'hFE644603;
    mem['h12D5] <= 32'hFE544783;
    mem['h12D6] <= 32'h00178793;
    mem['h12D7] <= 32'h00078693;
    mem['h12D8] <= 32'h00070513;
    mem['h12D9] <= 32'hA39FE0EF;
    mem['h12DA] <= 32'h00050793;
    mem['h12DB] <= 32'h00078663;
    mem['h12DC] <= 32'h00100793;
    mem['h12DD] <= 32'h0080006F;
    mem['h12DE] <= 32'h00000793;
    mem['h12DF] <= 32'h0FF7F713;
    mem['h12E0] <= 32'hFE544783;
    mem['h12E1] <= 32'h00F707B3;
    mem['h12E2] <= 32'hFEF402A3;
    mem['h12E3] <= 32'hFEB44783;
    mem['h12E4] <= 32'h02078A63;
    mem['h12E5] <= 32'hFE845703;
    mem['h12E6] <= 32'hFE744583;
    mem['h12E7] <= 32'hFE644783;
    mem['h12E8] <= 32'hFFF78793;
    mem['h12E9] <= 32'hFE544683;
    mem['h12EA] <= 32'h00078613;
    mem['h12EB] <= 32'h00070513;
    mem['h12EC] <= 32'h9EDFE0EF;
    mem['h12ED] <= 32'h00050793;
    mem['h12EE] <= 32'h00078663;
    mem['h12EF] <= 32'h00100793;
    mem['h12F0] <= 32'h0080006F;
    mem['h12F1] <= 32'h00000793;
    mem['h12F2] <= 32'h0FF7F793;
    mem['h12F3] <= 32'hFE644703;
    mem['h12F4] <= 32'h40F707B3;
    mem['h12F5] <= 32'hFEF40323;
    mem['h12F6] <= 32'hFED44783;
    mem['h12F7] <= 32'h04078C63;
    mem['h12F8] <= 32'hFE144783;
    mem['h12F9] <= 32'h02078A63;
    mem['h12FA] <= 32'hFE845703;
    mem['h12FB] <= 32'hFE744783;
    mem['h12FC] <= 32'h00178793;
    mem['h12FD] <= 32'hFE644603;
    mem['h12FE] <= 32'hFE544683;
    mem['h12FF] <= 32'h00078593;
    mem['h1300] <= 32'h00070513;
    mem['h1301] <= 32'h999FE0EF;
    mem['h1302] <= 32'h00050793;
    mem['h1303] <= 32'h00078663;
    mem['h1304] <= 32'h00100793;
    mem['h1305] <= 32'h0080006F;
    mem['h1306] <= 32'h00000793;
    mem['h1307] <= 32'h0FF7F713;
    mem['h1308] <= 32'hFE744783;
    mem['h1309] <= 32'h00F707B3;
    mem['h130A] <= 32'hFEF403A3;
    mem['h130B] <= 32'hFE0400A3;
    mem['h130C] <= 32'h00C0006F;
    mem['h130D] <= 32'h00100793;
    mem['h130E] <= 32'hFEF400A3;
    mem['h130F] <= 32'hFA144783;
    mem['h1310] <= 32'h3A078663;
    mem['h1311] <= 32'hFE0401A3;
    mem['h1312] <= 32'hFDE45783;
    mem['h1313] <= 32'h00178793;
    mem['h1314] <= 32'hFCF41F23;
    mem['h1315] <= 32'hFDE45703;
    mem['h1316] <= 32'h03200793;
    mem['h1317] <= 32'h02F777B3;
    mem['h1318] <= 32'h01079793;
    mem['h1319] <= 32'h0107D793;
    mem['h131A] <= 32'h00079E63;
    mem['h131B] <= 32'hFE444703;
    mem['h131C] <= 32'h00900793;
    mem['h131D] <= 32'h00E7F863;
    mem['h131E] <= 32'hFE444783;
    mem['h131F] <= 32'hFFF78793;
    mem['h1320] <= 32'hFEF40223;
    mem['h1321] <= 32'hFE845703;
    mem['h1322] <= 32'hFE744583;
    mem['h1323] <= 32'hFE644783;
    mem['h1324] <= 32'h00178793;
    mem['h1325] <= 32'hFE544683;
    mem['h1326] <= 32'h00078613;
    mem['h1327] <= 32'h00070513;
    mem['h1328] <= 32'h8FDFE0EF;
    mem['h1329] <= 32'h00050793;
    mem['h132A] <= 32'h00078E63;
    mem['h132B] <= 32'hFD644783;
    mem['h132C] <= 32'h00079A63;
    mem['h132D] <= 32'hFE644783;
    mem['h132E] <= 32'h00178793;
    mem['h132F] <= 32'hFEF40323;
    mem['h1330] <= 32'h32C0006F;
    mem['h1331] <= 32'hFE845703;
    mem['h1332] <= 32'hFE744583;
    mem['h1333] <= 32'hFE644783;
    mem['h1334] <= 32'hFFF78793;
    mem['h1335] <= 32'hFE544683;
    mem['h1336] <= 32'h00078613;
    mem['h1337] <= 32'h00070513;
    mem['h1338] <= 32'h8BDFE0EF;
    mem['h1339] <= 32'h00050793;
    mem['h133A] <= 32'h00078E63;
    mem['h133B] <= 32'hFD644783;
    mem['h133C] <= 32'h00078A63;
    mem['h133D] <= 32'hFE644783;
    mem['h133E] <= 32'hFFF78793;
    mem['h133F] <= 32'hFEF40323;
    mem['h1340] <= 32'h2EC0006F;
    mem['h1341] <= 32'hFC042623;
    mem['h1342] <= 32'h0B00006F;
    mem['h1343] <= 32'hFC042423;
    mem['h1344] <= 32'h0900006F;
    mem['h1345] <= 32'hFE845483;
    mem['h1346] <= 32'hFE744783;
    mem['h1347] <= 32'h00078613;
    mem['h1348] <= 32'hFC842583;
    mem['h1349] <= 32'hFCC42503;
    mem['h134A] <= 32'hF88FE0EF;
    mem['h134B] <= 32'h00050693;
    mem['h134C] <= 32'h00000713;
    mem['h134D] <= 32'h00449793;
    mem['h134E] <= 32'h00F707B3;
    mem['h134F] <= 32'h00D787B3;
    mem['h1350] <= 32'h0007C783;
    mem['h1351] <= 32'h04078863;
    mem['h1352] <= 32'hFE845783;
    mem['h1353] <= 32'h0FF7F693;
    mem['h1354] <= 32'hFE544703;
    mem['h1355] <= 32'hFC842783;
    mem['h1356] <= 32'h00F70733;
    mem['h1357] <= 32'h00070793;
    mem['h1358] <= 32'h00279793;
    mem['h1359] <= 32'h00E787B3;
    mem['h135A] <= 32'h00379793;
    mem['h135B] <= 32'h00078613;
    mem['h135C] <= 32'hFE644703;
    mem['h135D] <= 32'hFCC42783;
    mem['h135E] <= 32'h00F707B3;
    mem['h135F] <= 32'h00F607B3;
    mem['h1360] <= 32'h00168713;
    mem['h1361] <= 32'h0FF77713;
    mem['h1362] <= 32'h07C00693;
    mem['h1363] <= 32'h00F687B3;
    mem['h1364] <= 32'h00E78023;
    mem['h1365] <= 32'hFC842783;
    mem['h1366] <= 32'h00178793;
    mem['h1367] <= 32'hFCF42423;
    mem['h1368] <= 32'hFC842703;
    mem['h1369] <= 32'h00300793;
    mem['h136A] <= 32'hF6E7D6E3;
    mem['h136B] <= 32'hFCC42783;
    mem['h136C] <= 32'h00178793;
    mem['h136D] <= 32'hFCF42623;
    mem['h136E] <= 32'hFCC42703;
    mem['h136F] <= 32'h00300793;
    mem['h1370] <= 32'hF4E7D6E3;
    mem['h1371] <= 32'hFC042223;
    mem['h1372] <= 32'h13C0006F;
    mem['h1373] <= 32'h00100793;
    mem['h1374] <= 32'hFCF401A3;
    mem['h1375] <= 32'h00100793;
    mem['h1376] <= 32'hFAF42E23;
    mem['h1377] <= 32'h0840006F;
    mem['h1378] <= 32'hFE644703;
    mem['h1379] <= 32'hFC442783;
    mem['h137A] <= 32'h00F706B3;
    mem['h137B] <= 32'hFBC42703;
    mem['h137C] <= 32'h00070793;
    mem['h137D] <= 32'h00279793;
    mem['h137E] <= 32'h00E787B3;
    mem['h137F] <= 32'h00379793;
    mem['h1380] <= 32'h00F687B3;
    mem['h1381] <= 32'h07C00713;
    mem['h1382] <= 32'h00F707B3;
    mem['h1383] <= 32'h0007C783;
    mem['h1384] <= 32'h02078E63;
    mem['h1385] <= 32'hFE644703;
    mem['h1386] <= 32'hFC442783;
    mem['h1387] <= 32'h00F706B3;
    mem['h1388] <= 32'hFBC42703;
    mem['h1389] <= 32'h00070793;
    mem['h138A] <= 32'h00279793;
    mem['h138B] <= 32'h00E787B3;
    mem['h138C] <= 32'h00379793;
    mem['h138D] <= 32'h00F687B3;
    mem['h138E] <= 32'h07C00713;
    mem['h138F] <= 32'h00F707B3;
    mem['h1390] <= 32'h0007C703;
    mem['h1391] <= 32'h00900793;
    mem['h1392] <= 32'h00F71663;
    mem['h1393] <= 32'hFC0401A3;
    mem['h1394] <= 32'h01C0006F;
    mem['h1395] <= 32'hFBC42783;
    mem['h1396] <= 32'h00178793;
    mem['h1397] <= 32'hFAF42E23;
    mem['h1398] <= 32'hFBC42703;
    mem['h1399] <= 32'h01600793;
    mem['h139A] <= 32'hF6E7DCE3;
    mem['h139B] <= 32'hFC344783;
    mem['h139C] <= 32'h08078463;
    mem['h139D] <= 32'h00100793;
    mem['h139E] <= 32'hFAF42C23;
    mem['h139F] <= 32'h0400006F;
    mem['h13A0] <= 32'hFE644703;
    mem['h13A1] <= 32'hFC442783;
    mem['h13A2] <= 32'h00F706B3;
    mem['h13A3] <= 32'hFB842703;
    mem['h13A4] <= 32'h00070793;
    mem['h13A5] <= 32'h00279793;
    mem['h13A6] <= 32'h00E787B3;
    mem['h13A7] <= 32'h00379793;
    mem['h13A8] <= 32'h00F687B3;
    mem['h13A9] <= 32'h07C00713;
    mem['h13AA] <= 32'h00F707B3;
    mem['h13AB] <= 32'h00078023;
    mem['h13AC] <= 32'hFB842783;
    mem['h13AD] <= 32'h00178793;
    mem['h13AE] <= 32'hFAF42C23;
    mem['h13AF] <= 32'hFB842703;
    mem['h13B0] <= 32'h01600793;
    mem['h13B1] <= 32'hFAE7DEE3;
    mem['h13B2] <= 32'hFC442783;
    mem['h13B3] <= 32'h0FF7F693;
    mem['h13B4] <= 32'hFDB44783;
    mem['h13B5] <= 32'hFE644703;
    mem['h13B6] <= 32'h00E68733;
    mem['h13B7] <= 32'h0FF77713;
    mem['h13B8] <= 32'hFF040693;
    mem['h13B9] <= 32'h00F687B3;
    mem['h13BA] <= 32'hFAE78623;
    mem['h13BB] <= 32'hFDB44783;
    mem['h13BC] <= 32'h00178793;
    mem['h13BD] <= 32'hFCF40DA3;
    mem['h13BE] <= 32'hFC442783;
    mem['h13BF] <= 32'h00178793;
    mem['h13C0] <= 32'hFCF42223;
    mem['h13C1] <= 32'hFC442703;
    mem['h13C2] <= 32'h00300793;
    mem['h13C3] <= 32'hECE7D0E3;
    mem['h13C4] <= 32'hFD644783;
    mem['h13C5] <= 32'hFCF40C23;
    mem['h13C6] <= 32'hFDC45783;
    mem['h13C7] <= 32'h00178793;
    mem['h13C8] <= 32'hFCF41E23;
    mem['h13C9] <= 32'hFDB44783;
    mem['h13CA] <= 32'h02078263;
    mem['h13CB] <= 32'hFDB44783;
    mem['h13CC] <= 32'h01400713;
    mem['h13CD] <= 32'h00F717B3;
    mem['h13CE] <= 32'h01079713;
    mem['h13CF] <= 32'h01075713;
    mem['h13D0] <= 32'hFDC45783;
    mem['h13D1] <= 32'h00F707B3;
    mem['h13D2] <= 32'hFCF41E23;
    mem['h13D3] <= 32'h00100793;
    mem['h13D4] <= 32'hFCF40BA3;
    mem['h13D5] <= 32'h01300593;
    mem['h13D6] <= 32'h00200513;
    mem['h13D7] <= 32'hE40FF0EF;
    mem['h13D8] <= 32'h00050793;
    mem['h13D9] <= 32'hFEF402A3;
    mem['h13DA] <= 32'hE00FF0EF;
    mem['h13DB] <= 32'h00050793;
    mem['h13DC] <= 32'hFCF40B23;
    mem['h13DD] <= 32'hFD644783;
    mem['h13DE] <= 32'h00079A63;
    mem['h13DF] <= 32'h00300793;
    mem['h13E0] <= 32'hFEF403A3;
    mem['h13E1] <= 32'hFE040323;
    mem['h13E2] <= 32'h0140006F;
    mem['h13E3] <= 32'h00300793;
    mem['h13E4] <= 32'hFEF403A3;
    mem['h13E5] <= 32'h02400793;
    mem['h13E6] <= 32'hFEF40323;
    mem['h13E7] <= 32'hFDE45703;
    mem['h13E8] <= 32'h00700793;
    mem['h13E9] <= 32'h02F777B3;
    mem['h13EA] <= 32'hFEF41423;
    mem['h13EB] <= 32'hFE845783;
    mem['h13EC] <= 32'hFE744703;
    mem['h13ED] <= 32'hFE644603;
    mem['h13EE] <= 32'hFE544683;
    mem['h13EF] <= 32'h00070593;
    mem['h13F0] <= 32'h00078513;
    mem['h13F1] <= 32'hDD8FE0EF;
    mem['h13F2] <= 32'h00050793;
    mem['h13F3] <= 32'h00F037B3;
    mem['h13F4] <= 32'h0FF7F793;
    mem['h13F5] <= 32'h0017C793;
    mem['h13F6] <= 32'h0FF7F793;
    mem['h13F7] <= 32'hFCF40D23;
    mem['h13F8] <= 32'hFDA44783;
    mem['h13F9] <= 32'h0017F793;
    mem['h13FA] <= 32'hFCF40D23;
    mem['h13FB] <= 32'hFD744783;
    mem['h13FC] <= 32'h00078E63;
    mem['h13FD] <= 32'hFC040BA3;
    mem['h13FE] <= 32'hFDC45783;
    mem['h13FF] <= 32'h01800613;
    mem['h1400] <= 32'h01600593;
    mem['h1401] <= 32'h00078513;
    mem['h1402] <= 32'hE1DFE0EF;
    mem['h1403] <= 32'hFA042A23;
    mem['h1404] <= 32'h0900006F;
    mem['h1405] <= 32'hFA042823;
    mem['h1406] <= 32'h0700006F;
    mem['h1407] <= 32'hFB442703;
    mem['h1408] <= 32'h00070793;
    mem['h1409] <= 32'h00279793;
    mem['h140A] <= 32'h00E787B3;
    mem['h140B] <= 32'h00379793;
    mem['h140C] <= 32'h00078713;
    mem['h140D] <= 32'hFB042783;
    mem['h140E] <= 32'h00F707B3;
    mem['h140F] <= 32'h07C00713;
    mem['h1410] <= 32'h00F707B3;
    mem['h1411] <= 32'h0007C683;
    mem['h1412] <= 32'hFB442703;
    mem['h1413] <= 32'h00070793;
    mem['h1414] <= 32'h00279793;
    mem['h1415] <= 32'h00E787B3;
    mem['h1416] <= 32'h00379793;
    mem['h1417] <= 32'h00078713;
    mem['h1418] <= 32'hFB042783;
    mem['h1419] <= 32'h00F707B3;
    mem['h141A] <= 32'h00279713;
    mem['h141B] <= 32'h052007B7;
    mem['h141C] <= 32'h00F707B3;
    mem['h141D] <= 32'h00068713;
    mem['h141E] <= 32'h00E7A023;
    mem['h141F] <= 32'hFB042783;
    mem['h1420] <= 32'h00178793;
    mem['h1421] <= 32'hFAF42823;
    mem['h1422] <= 32'hFB042703;
    mem['h1423] <= 32'h02700793;
    mem['h1424] <= 32'hF8E7D6E3;
    mem['h1425] <= 32'hFB442783;
    mem['h1426] <= 32'h00178793;
    mem['h1427] <= 32'hFAF42A23;
    mem['h1428] <= 32'hFB442703;
    mem['h1429] <= 32'h01D00793;
    mem['h142A] <= 32'hF6E7D6E3;
    mem['h142B] <= 32'hFA042623;
    mem['h142C] <= 32'h0B00006F;
    mem['h142D] <= 32'hFA042423;
    mem['h142E] <= 32'h0900006F;
    mem['h142F] <= 32'hFE845483;
    mem['h1430] <= 32'hFE744783;
    mem['h1431] <= 32'h00078613;
    mem['h1432] <= 32'hFA842583;
    mem['h1433] <= 32'hFAC42503;
    mem['h1434] <= 32'hBE0FE0EF;
    mem['h1435] <= 32'h00050693;
    mem['h1436] <= 32'h00000713;
    mem['h1437] <= 32'h00449793;
    mem['h1438] <= 32'h00F707B3;
    mem['h1439] <= 32'h00D787B3;
    mem['h143A] <= 32'h0007C783;
    mem['h143B] <= 32'h04078863;
    mem['h143C] <= 32'hFE845783;
    mem['h143D] <= 32'h00178693;
    mem['h143E] <= 32'hFE544703;
    mem['h143F] <= 32'hFA842783;
    mem['h1440] <= 32'h00F70733;
    mem['h1441] <= 32'h00070793;
    mem['h1442] <= 32'h00279793;
    mem['h1443] <= 32'h00E787B3;
    mem['h1444] <= 32'h00379793;
    mem['h1445] <= 32'h00078613;
    mem['h1446] <= 32'hFE644703;
    mem['h1447] <= 32'hFAC42783;
    mem['h1448] <= 32'h00F707B3;
    mem['h1449] <= 32'h00F607B3;
    mem['h144A] <= 32'h00279713;
    mem['h144B] <= 32'h052007B7;
    mem['h144C] <= 32'h00F707B3;
    mem['h144D] <= 32'h00068713;
    mem['h144E] <= 32'h00E7A023;
    mem['h144F] <= 32'hFA842783;
    mem['h1450] <= 32'h00178793;
    mem['h1451] <= 32'hFAF42423;
    mem['h1452] <= 32'hFA842703;
    mem['h1453] <= 32'h00300793;
    mem['h1454] <= 32'hF6E7D6E3;
    mem['h1455] <= 32'hFAC42783;
    mem['h1456] <= 32'h00178793;
    mem['h1457] <= 32'hFAF42623;
    mem['h1458] <= 32'hFAC42703;
    mem['h1459] <= 32'h00300793;
    mem['h145A] <= 32'hF4E7D6E3;
    mem['h145B] <= 32'hFDB44783;
    mem['h145C] <= 32'h1A078A63;
    mem['h145D] <= 32'hFD844783;
    mem['h145E] <= 32'h0C079663;
    mem['h145F] <= 32'hFA0403A3;
    mem['h1460] <= 32'h0B40006F;
    mem['h1461] <= 32'hFA744783;
    mem['h1462] <= 32'hFF040713;
    mem['h1463] <= 32'h00F707B3;
    mem['h1464] <= 32'hFAC7C783;
    mem['h1465] <= 32'hFAF40323;
    mem['h1466] <= 32'h0880006F;
    mem['h1467] <= 32'h00100793;
    mem['h1468] <= 32'hFAF402A3;
    mem['h1469] <= 32'h0640006F;
    mem['h146A] <= 32'hFA644783;
    mem['h146B] <= 32'hFFF78693;
    mem['h146C] <= 32'hFA544703;
    mem['h146D] <= 32'h00070793;
    mem['h146E] <= 32'h00279793;
    mem['h146F] <= 32'h00E787B3;
    mem['h1470] <= 32'h00379793;
    mem['h1471] <= 32'h00F686B3;
    mem['h1472] <= 32'hFA644603;
    mem['h1473] <= 32'hFA544703;
    mem['h1474] <= 32'h00070793;
    mem['h1475] <= 32'h00279793;
    mem['h1476] <= 32'h00E787B3;
    mem['h1477] <= 32'h00379793;
    mem['h1478] <= 32'h00F607B3;
    mem['h1479] <= 32'h07C00713;
    mem['h147A] <= 32'h00D70733;
    mem['h147B] <= 32'h00074703;
    mem['h147C] <= 32'h07C00693;
    mem['h147D] <= 32'h00F687B3;
    mem['h147E] <= 32'h00E78023;
    mem['h147F] <= 32'hFA544783;
    mem['h1480] <= 32'h00178793;
    mem['h1481] <= 32'hFAF402A3;
    mem['h1482] <= 32'hFA544703;
    mem['h1483] <= 32'h01600793;
    mem['h1484] <= 32'hF8E7FCE3;
    mem['h1485] <= 32'hFA644783;
    mem['h1486] <= 32'hFFF78793;
    mem['h1487] <= 32'hFAF40323;
    mem['h1488] <= 32'hFA644783;
    mem['h1489] <= 32'hF6079CE3;
    mem['h148A] <= 32'hFA744783;
    mem['h148B] <= 32'h00178793;
    mem['h148C] <= 32'hFAF403A3;
    mem['h148D] <= 32'hFA744703;
    mem['h148E] <= 32'hFDB44783;
    mem['h148F] <= 32'hF4F764E3;
    mem['h1490] <= 32'h0D00006F;
    mem['h1491] <= 32'hFDB44783;
    mem['h1492] <= 32'hFAF40223;
    mem['h1493] <= 32'h0BC0006F;
    mem['h1494] <= 32'hFA444783;
    mem['h1495] <= 32'hFFF78793;
    mem['h1496] <= 32'hFF040713;
    mem['h1497] <= 32'h00F707B3;
    mem['h1498] <= 32'hFAC7C783;
    mem['h1499] <= 32'hFAF401A3;
    mem['h149A] <= 32'h0880006F;
    mem['h149B] <= 32'h00100793;
    mem['h149C] <= 32'hFAF40123;
    mem['h149D] <= 32'h0640006F;
    mem['h149E] <= 32'hFA344783;
    mem['h149F] <= 32'h00178693;
    mem['h14A0] <= 32'hFA244703;
    mem['h14A1] <= 32'h00070793;
    mem['h14A2] <= 32'h00279793;
    mem['h14A3] <= 32'h00E787B3;
    mem['h14A4] <= 32'h00379793;
    mem['h14A5] <= 32'h00F686B3;
    mem['h14A6] <= 32'hFA344603;
    mem['h14A7] <= 32'hFA244703;
    mem['h14A8] <= 32'h00070793;
    mem['h14A9] <= 32'h00279793;
    mem['h14AA] <= 32'h00E787B3;
    mem['h14AB] <= 32'h00379793;
    mem['h14AC] <= 32'h00F607B3;
    mem['h14AD] <= 32'h07C00713;
    mem['h14AE] <= 32'h00D70733;
    mem['h14AF] <= 32'h00074703;
    mem['h14B0] <= 32'h07C00693;
    mem['h14B1] <= 32'h00F687B3;
    mem['h14B2] <= 32'h00E78023;
    mem['h14B3] <= 32'hFA244783;
    mem['h14B4] <= 32'h00178793;
    mem['h14B5] <= 32'hFAF40123;
    mem['h14B6] <= 32'hFA244703;
    mem['h14B7] <= 32'h01600793;
    mem['h14B8] <= 32'hF8E7FCE3;
    mem['h14B9] <= 32'hFA344783;
    mem['h14BA] <= 32'h00178793;
    mem['h14BB] <= 32'hFAF401A3;
    mem['h14BC] <= 32'hFA344703;
    mem['h14BD] <= 32'h02600793;
    mem['h14BE] <= 32'hF6E7FAE3;
    mem['h14BF] <= 32'hFA444783;
    mem['h14C0] <= 32'hFFF78793;
    mem['h14C1] <= 32'hFAF40223;
    mem['h14C2] <= 32'hFA444783;
    mem['h14C3] <= 32'hF40792E3;
    mem['h14C4] <= 32'hF8040E23;
    mem['h14C5] <= 32'hF8040EA3;
    mem['h14C6] <= 32'hF8040F23;
    mem['h14C7] <= 32'hF8040FA3;
    mem['h14C8] <= 32'hFC040DA3;
    mem['h14C9] <= 32'hFE0407A3;
    mem['h14CA] <= 32'hFE040723;
    mem['h14CB] <= 32'hFE0406A3;
    mem['h14CC] <= 32'hFE040623;
    mem['h14CD] <= 32'hFE0405A3;
    mem['h14CE] <= 32'hBF8FF06F;
    mem['h14CF] <= 32'hFE010113;
    mem['h14D0] <= 32'h00112E23;
    mem['h14D1] <= 32'h00812C23;
    mem['h14D2] <= 32'h02010413;
    mem['h14D3] <= 32'h00050793;
    mem['h14D4] <= 32'hFEF407A3;
    mem['h14D5] <= 32'hFEF44703;
    mem['h14D6] <= 32'h00A00793;
    mem['h14D7] <= 32'h00F71663;
    mem['h14D8] <= 32'h00D00513;
    mem['h14D9] <= 32'hFD9FF0EF;
    mem['h14DA] <= 32'h020007B7;
    mem['h14DB] <= 32'h00878793;
    mem['h14DC] <= 32'hFEF44703;
    mem['h14DD] <= 32'h00E7A023;
    mem['h14DE] <= 32'h00000013;
    mem['h14DF] <= 32'h01C12083;
    mem['h14E0] <= 32'h01812403;
    mem['h14E1] <= 32'h02010113;
    mem['h14E2] <= 32'h00008067;
    mem['h14E3] <= 32'hFE010113;
    mem['h14E4] <= 32'h00112E23;
    mem['h14E5] <= 32'h00812C23;
    mem['h14E6] <= 32'h02010413;
    mem['h14E7] <= 32'hFEA42623;
    mem['h14E8] <= 32'h01C0006F;
    mem['h14E9] <= 32'hFEC42783;
    mem['h14EA] <= 32'h00178713;
    mem['h14EB] <= 32'hFEE42623;
    mem['h14EC] <= 32'h0007C783;
    mem['h14ED] <= 32'h00078513;
    mem['h14EE] <= 32'hF85FF0EF;
    mem['h14EF] <= 32'hFEC42783;
    mem['h14F0] <= 32'h0007C783;
    mem['h14F1] <= 32'hFE0790E3;
    mem['h14F2] <= 32'h00000013;
    mem['h14F3] <= 32'h00000013;
    mem['h14F4] <= 32'h01C12083;
    mem['h14F5] <= 32'h01812403;
    mem['h14F6] <= 32'h02010113;
    mem['h14F7] <= 32'h00008067;
    mem['h14F8] <= 32'hFD010113;
    mem['h14F9] <= 32'h02812623;
    mem['h14FA] <= 32'h03010413;
    mem['h14FB] <= 32'hFCA42E23;
    mem['h14FC] <= 32'hFCB42C23;
    mem['h14FD] <= 32'hFD842783;
    mem['h14FE] <= 32'hFFF78793;
    mem['h14FF] <= 32'h00279793;
    mem['h1500] <= 32'hFEF42623;
    mem['h1501] <= 32'h03C0006F;
    mem['h1502] <= 32'hFEC42783;
    mem['h1503] <= 32'hFDC42703;
    mem['h1504] <= 32'h00F757B3;
    mem['h1505] <= 32'h00F7F793;
    mem['h1506] <= 32'h00105737;
    mem['h1507] <= 32'h4F070713;
    mem['h1508] <= 32'h00F707B3;
    mem['h1509] <= 32'h0007C703;
    mem['h150A] <= 32'h020007B7;
    mem['h150B] <= 32'h00878793;
    mem['h150C] <= 32'h00E7A023;
    mem['h150D] <= 32'hFEC42783;
    mem['h150E] <= 32'hFFC78793;
    mem['h150F] <= 32'hFEF42623;
    mem['h1510] <= 32'hFEC42783;
    mem['h1511] <= 32'hFC07D2E3;
    mem['h1512] <= 32'h00000013;
    mem['h1513] <= 32'h00000013;
    mem['h1514] <= 32'h02C12403;
    mem['h1515] <= 32'h03010113;
    mem['h1516] <= 32'h00008067;
    mem['h1517] <= 32'h00103738;
    mem['h1518] <= 32'h001037D4;
    mem['h1519] <= 32'h00103858;
    mem['h151A] <= 32'h00103924;
    mem['h151B] <= 32'h001039C4;
    mem['h151C] <= 32'h00103A64;
    mem['h151D] <= 32'h00103B30;
    mem['h151E] <= 32'h00103BEC;
    mem['h151F] <= 32'h00103C6C;
    mem['h1520] <= 32'h00103D18;
    mem['h1521] <= 32'h6C65645F;
    mem['h1522] <= 32'h63207961;
    mem['h1523] <= 32'h656C6C61;
    mem['h1524] <= 32'h00000064;
    mem['h1525] <= 32'h72746554;
    mem['h1526] <= 32'h72615369;
    mem['h1527] <= 32'h0A216A61;
    mem['h1528] <= 32'h00000000;
    mem['h1529] <= 32'h54545542;
    mem['h152A] <= 32'h555F4E4F;
    mem['h152B] <= 32'h00000A50;
    mem['h152C] <= 32'h54545542;
    mem['h152D] <= 32'h445F4E4F;
    mem['h152E] <= 32'h0A4E574F;
    mem['h152F] <= 32'h00000000;
    mem['h1530] <= 32'h54545542;
    mem['h1531] <= 32'h525F4E4F;
    mem['h1532] <= 32'h54484749;
    mem['h1533] <= 32'h0000000A;
    mem['h1534] <= 32'h54545542;
    mem['h1535] <= 32'h4C5F4E4F;
    mem['h1536] <= 32'h0A544645;
    mem['h1537] <= 32'h00000000;
    mem['h1538] <= 32'h54545542;
    mem['h1539] <= 32'h435F4E4F;
    mem['h153A] <= 32'h45544E45;
    mem['h153B] <= 32'h00000A52;
    mem['h153C] <= 32'h33323130;
    mem['h153D] <= 32'h37363534;
    mem['h153E] <= 32'h42413938;
    mem['h153F] <= 32'h46454443;
    mem['h1540] <= 32'h00000000;
    mem['h1541] <= 32'h01010101;
    mem['h1542] <= 32'h00000000;
    mem['h1543] <= 32'h00000000;
    mem['h1544] <= 32'h00000000;
    mem['h1545] <= 32'h00010000;
    mem['h1546] <= 32'h00010100;
    mem['h1547] <= 32'h00010000;
    mem['h1548] <= 32'h00000000;
    mem['h1549] <= 32'h00000000;
    mem['h154A] <= 32'h00010100;
    mem['h154B] <= 32'h00010100;
    mem['h154C] <= 32'h00000000;
    mem['h154D] <= 32'h00010000;
    mem['h154E] <= 32'h00010100;
    mem['h154F] <= 32'h00000100;
    mem['h1550] <= 32'h00000000;
    mem['h1551] <= 32'h00000100;
    mem['h1552] <= 32'h00010100;
    mem['h1553] <= 32'h00010000;
    mem['h1554] <= 32'h00000000;
    mem['h1555] <= 32'h00000100;
    mem['h1556] <= 32'h00000100;
    mem['h1557] <= 32'h00010100;
    mem['h1558] <= 32'h00000000;
    mem['h1559] <= 32'h00010000;
    mem['h155A] <= 32'h00010000;
    mem['h155B] <= 32'h00010100;
    mem['h155C] <= 32'h00000000;
    mem['h155D] <= 32'h000009C4;
    mem['h155E] <= 32'h075BCD15;
    mem['h155F] <= 32'h075BCD15;

  end

  always @(posedge clk) mem_data <= mem[mem_addr];

  // ============================================================================

  reg o_ready;

  always @(posedge clk or negedge rstn)
    if (!rstn) o_ready <= 1'd0;
    else o_ready <= valid && ((addr & MEM_ADDR_MASK) != 0);

  // Output connectins
  assign ready    = o_ready;
  assign rdata    = mem_data;
  assign mem_addr = addr[MEM_SIZE_BITS+1:2];

  always @(posedge clk) begin    
    if (wen) mem[waddr] <= wdata;				
  end

endmodule
