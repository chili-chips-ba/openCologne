//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 May 2024)
//  Compile Time: 1970-01-01 00:59:59
//  Program Run:  2024-07-11 21:42:09
//  Program Call: p_r +sp -i /home/user/FPGA/Boards/GateMate/gatemate_ila/net/ila_top_synth24-07-11_21-41-30.v -o /home/user/FPGA/Boards/GateMate/gatemate_ila/p_r_out/ila_top_24-07-11_21-41-30 -sp -cCP +uCIO -ccf /home/user/FPGA/Boards/GateMate/gatemate_ila/src/ILA_top.ccf 
//  File Type:    Verilog

// Gatecount:    305
module ila_top_24-07-11_21-41-30 (clk , i_mosi_ILA , i_sclk_ILA , i_ss_ILA ,
       led , o_miso_ILA 
       ) ;

input  clk;
input  i_mosi_ILA;
input  i_sclk_ILA;
input  i_ss_ILA;

output led;
output o_miso_ILA;



wire clk;
wire led;
wire na1_1;
wire na1_1_i;
wire na2_2;
wire na4_1;
wire na5_1;
wire na6_1;
wire na6_1_i;
wire na6_2;
wire na6_2_i;
wire na8_1;
wire na8_1_i;
wire na9_1;
wire na9_1_i;
wire na9_2;
wire na9_2_i;
wire na10_1;
wire na10_1_i;
wire na11_1;
wire na11_1_i;
wire na12_1;
wire na12_1_i;
wire na13_1;
wire na14_1;
wire na14_1_i;
wire na14_2;
wire na14_2_i;
wire na15_1;
wire na15_1_i;
wire na18_2;
wire na18_2_i;
wire na19_1;
wire na19_1_i;
wire na19_2;
wire na19_2_i;
wire na20_1;
wire na20_1_i;
wire na20_2;
wire na20_2_i;
wire na22_1;
wire na22_1_i;
wire na22_2;
wire na22_2_i;
wire na23_1;
wire na23_1_i;
wire na23_2;
wire na23_2_i;
wire na24_1;
wire na24_1_i;
wire na26_1;
wire na26_1_i;
wire na26_2;
wire na26_2_i;
wire na27_1;
wire na27_1_i;
wire na27_2;
wire na27_2_i;
wire na28_1;
wire na28_1_i;
wire na28_2;
wire na28_2_i;
wire na29_2;
wire na29_2_i;
wire na30_1;
wire na30_1_i;
wire na30_2;
wire na30_2_i;
wire na31_1;
wire na31_1_i;
wire na31_2;
wire na31_2_i;
wire na33_1;
wire na33_1_i;
wire na33_2;
wire na33_2_i;
wire na35_1;
wire na35_1_i;
wire na36_1;
wire na36_1_i;
wire na37_2;
wire na39_1;
wire na39_1_i;
wire na39_2;
wire na39_2_i;
wire na40_2;
wire na40_2_i;
wire na41_1;
wire na42_1;
wire na42_1_i;
wire na43_2;
wire na43_2_i;
wire na44_1;
wire na44_1_i;
wire na45_1;
wire na45_1_i;
wire na46_2;
wire na46_2_i;
wire na47_1;
wire na47_1_i;
wire na48_2;
wire na48_2_i;
wire na49_2;
wire na49_2_i;
wire na50_1;
wire na50_1_i;
wire na51_2;
wire na51_2_i;
wire na52_1;
wire na52_1_i;
wire na53_1;
wire na54_1;
wire na54_1_i;
wire na55_1;
wire na55_1_i;
wire na55_2;
wire na55_2_i;
wire na57_1;
wire na57_1_i;
wire na58_2;
wire na58_2_i;
wire na59_1;
wire na59_1_i;
wire na59_2;
wire na59_2_i;
wire na60_1;
wire na60_1_i;
wire na61_1;
wire na61_1_i;
wire na62_1;
wire na62_1_i;
wire na62_2;
wire na62_2_i;
wire na64_1;
wire na64_1_i;
wire na64_2;
wire na64_2_i;
wire na65_1;
wire na65_1_i;
wire na67_1;
wire na67_1_i;
wire na67_2;
wire na67_2_i;
wire na68_1;
wire na68_1_i;
wire na72_2;
wire na72_2_i;
wire na73_1;
wire na74_1;
wire na74_1_i;
wire na75_1;
wire na75_1_i;
wire na76_1;
wire na76_1_i;
wire na76_2;
wire na76_2_i;
wire na77_1;
wire na77_1_i;
wire na77_2;
wire na77_2_i;
wire na78_1;
wire na78_1_i;
wire na78_2;
wire na78_2_i;
wire na79_1;
wire na79_1_i;
wire na80_1;
wire na80_1_i;
wire na81_2;
wire na84_1;
wire na84_1_i;
wire na84_2;
wire na84_2_i;
wire na87_1;
wire na87_1_i;
wire na87_2;
wire na87_2_i;
wire na89_1;
wire na89_1_i;
wire na89_2;
wire na89_2_i;
wire na90_1;
wire na90_1_i;
wire na90_2;
wire na90_2_i;
wire na91_2;
wire na91_2_i;
wire na92_1;
wire na92_1_i;
wire na93_2;
wire na93_2_i;
wire na94_1;
wire na94_1_i;
wire na96_1;
wire na96_1_i;
wire na96_2;
wire na96_2_i;
wire na98_2;
wire na98_2_i;
wire na100_1;
wire na100_1_i;
wire na102_1;
wire na102_1_i;
wire na102_2;
wire na102_2_i;
wire na103_1;
wire na103_1_i;
wire na106_1;
wire na106_1_i;
wire na106_2;
wire na106_2_i;
wire na108_1;
wire na108_1_i;
wire na110_1;
wire na110_1_i;
wire na111_1;
wire na111_1_i;
wire na112_1;
wire na112_1_i;
wire na112_2;
wire na112_2_i;
wire na113_1;
wire na113_1_i;
wire na113_2;
wire na113_2_i;
wire na115_2;
wire na115_2_i;
wire na116_1;
wire na116_1_i;
wire na117_1;
wire na117_1_i;
wire na118_1;
wire na118_1_i;
wire na119_1;
wire na119_1_i;
wire na120_1;
wire na120_1_i;
wire na121_1;
wire na121_1_i;
wire na122_1;
wire na122_1_i;
wire na123_1;
wire na123_1_i;
wire na124_1;
wire na124_1_i;
wire na125_1;
wire na125_1_i;
wire na126_1;
wire na126_1_i;
wire na130_2;
wire na130_2_i;
wire na131_1;
wire na131_1_i;
wire na131_2;
wire na131_2_i;
wire na133_1;
wire na134_1;
wire na138_1;
wire na139_2;
wire na139_2_i;
wire na140_1;
wire na141_1;
wire na141_1_i;
wire na144_1;
wire na144_2;
wire na144_4;
wire na146_1;
wire na146_2;
wire na146_4;
wire na148_1;
wire na148_2;
wire na148_4;
wire na150_1;
wire na150_2;
wire na150_4;
wire na152_1;
wire na152_2;
wire na152_4;
wire na153_1;
wire na153_2;
wire na153_4;
wire na155_1;
wire na155_2;
wire na155_4;
wire na157_1;
wire na157_2;
wire na160_1;
wire na160_2;
wire na160_4;
wire na162_1;
wire na162_2;
wire na162_4;
wire na164_1;
wire na164_2;
wire na164_4;
wire na166_1;
wire na166_2;
wire na166_4;
wire na167_1;
wire na167_4;
wire na168_1;
wire na168_2;
wire na168_4;
wire na170_1;
wire na170_2;
wire na170_4;
wire na172_1;
wire na172_2;
wire na172_4;
wire na174_1;
wire na174_2;
wire na176_1;
wire na176_4;
wire na177_1;
wire na177_2;
wire na177_4;
wire na179_1;
wire na179_2;
wire na179_4;
wire na181_1;
wire na181_2;
wire na181_4;
wire na183_1;
wire na183_2;
wire na185_1;
wire na185_4;
wire na186_1;
wire na186_2;
wire na186_4;
wire na188_1;
wire na188_2;
wire na188_4;
wire na190_1;
wire na190_2;
wire na190_4;
wire na192_1;
wire na192_2;
wire na194_1;
wire na194_4;
wire na195_1;
wire na195_2;
wire na195_4;
wire na197_1;
wire na197_2;
wire na197_4;
wire na199_1;
wire na199_2;
wire na199_4;
wire na201_1;
wire na201_2;
wire na205_1;
wire na205_2;
wire na247_2;
wire na247_2_i;
wire na248_1;
wire na248_1_i;
wire na315_2;
wire na315_2_i;
wire na332_1;
wire na333_1;
wire na334_1;
wire na335_1;
wire na336_1;
wire na339_3;
wire na339_4;
wire na339_5;
wire na339_6;
wire na340_3;
wire na340_4;
wire na340_5;
wire na340_6;
wire na342_1;
wire na343_2;
wire na344_1;
wire na344_4;
wire na345_1;
wire na346_1;
wire na347_1;
wire na348_1;
wire na348_2;
wire na349_1;
wire na350_2;
wire na351_1;
wire na352_1;
wire na353_1;
wire na354_1;
wire na355_1;
wire na356_1;
wire na357_1;
wire na358_1;
wire na358_9;
wire na359_1;
wire na360_2;
wire na361_1;
wire na362_2;
wire na363_2;
wire na364_1;
wire na364_9;
wire na365_2;
wire na366_1;
wire na366_9;
wire na367_2;
wire na368_1;
wire na369_1;
wire na370_1;
wire na371_2;
wire na372_1;
wire na373_1;
wire na374_1;
wire na375_1;
wire na376_2;
wire na377_1;
wire na378_1;
wire na379_1;
wire na380_1;
wire na380_9;
wire na381_1;
wire na382_1;
wire na383_1;
wire na384_1;
wire na385_2;
wire na386_1;
wire na387_1;
wire na387_9;
wire na388_1;
wire na389_1;
wire na390_2;
wire na391_1;
wire na392_1;
wire na392_9;
wire na393_1;
wire na394_2;
wire na395_1;
wire na396_1;
wire na397_1;
wire na397_9;
wire na398_2;
wire na399_1;
wire na399_9;
wire na400_2;
wire na401_2;
wire na402_1;
wire na403_2;
wire na404_2;
wire na405_1;
wire na405_9;
wire na406_2;
wire na407_1;
wire na407_9;
wire na408_2;
wire na409_1;
wire na409_9;
wire na410_2;
wire na411_1;
wire na411_9;
wire na412_2;
wire na413_1;
wire na413_9;
wire na414_2;
wire na415_1;
wire na415_9;
wire na416_2;
wire na417_1;
wire na417_9;
wire na418_2;
wire na419_1;
wire na419_9;
wire na420_2;
wire na421_1;
wire na421_9;
wire na422_2;
wire na423_1;
wire na423_9;
wire na424_2;
wire na425_1;
wire na425_9;
wire na426_2;
wire na427_1;
wire na427_9;
wire na428_2;
wire na429_1;
wire na429_9;
wire na430_2;
wire na431_1;
wire na431_9;
wire na432_2;
wire na433_1;
wire na433_9;
wire na434_2;
wire na435_1;
wire na435_9;
wire na436_2;
wire na437_1;
wire na437_9;
wire na438_2;
wire na439_1;
wire na439_9;
wire na440_2;
wire na441_1;
wire na441_9;
wire na442_2;
wire na443_1;
wire na443_9;
wire na444_2;
wire na445_1;
wire na445_9;
wire na446_2;
wire na447_1;
wire na447_9;
wire na448_2;
wire na449_1;
wire na449_9;
wire na450_2;
wire na451_1;
wire na451_9;
wire na452_2;
wire na453_1;
wire na453_9;
wire na454_2;
wire na455_1;
wire na455_9;
wire na456_2;
wire na457_1;
wire na458_2;
wire na459_1;
wire na460_2;
wire na461_1;
wire na462_2;
wire na463_2;
wire na464_2;
wire na465_2;
wire na466_2;
wire na467_2;
wire na468_2;
wire na469_2;
wire na470_2;
wire na471_2;
wire na472_2;
wire na473_2;
wire na474_2;
wire na475_2;
wire na476_2;
wire na477_2;
wire na478_2;
wire na479_2;
wire na480_2;
wire na481_2;
wire na482_2;
wire na483_2;
wire na484_2;
wire na485_2;
wire na486_2;
wire na487_2;
wire na488_2;
wire na489_2;
wire na490_2;
wire na491_2;
wire na492_2;
wire na493_2;
wire na494_2;
wire na495_2;
wire na496_2;
wire na497_2;
wire na498_2;
wire na499_2;
wire na500_2;
wire na501_2;
wire i_ss_ILA;
wire na341_96;
wire na341_97;
wire na341_98;
wire na341_99;
wire na360_10;
wire na362_10;
wire na365_10;
wire na376_10;
wire na385_10;
wire na390_10;
wire na394_10;
wire na398_10;
wire na400_10;
wire na403_10;
wire na404_10;
wire na406_10;
wire na408_10;
wire na410_10;
wire na412_10;
wire na414_10;
wire na416_10;
wire na418_10;
wire na420_10;
wire na422_10;
wire na424_10;
wire na426_10;
wire na428_10;
wire na430_10;
wire na432_10;
wire na434_10;
wire na436_10;
wire na438_10;
wire na440_10;
wire na442_10;
wire na444_10;
wire na446_10;
wire na448_10;
wire na450_10;
wire na452_10;
wire na454_10;
wire na456_10;
wire na341_100;
wire i_mosi_ILA;
wire i_sclk_ILA;
wire o_miso_ILA;

// C_ORAND/D///      x17y38     80'h00_FD00_00_0000_0888_3FCE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1_1 ( .OUT(na1_1_i), .IN1(na2_2), .IN2(na12_1), .IN3(1'b0), .IN4(na343_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0), .IN8(~na336_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1_2 ( .OUT(na1_1), .CLK(~na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1_1_i) );
// C_///AND/      x17y37     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2_4 ( .OUT(na2_2), .IN1(na14_1), .IN2(1'b1), .IN3(na465_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x19y40     80'h00_0018_00_0000_0C88_8CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4_1 ( .OUT(na4_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na26_2), .IN7(na39_2), .IN8(na47_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x22y42     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a5_1 ( .OUT(na5_1), .IN1(1'b1), .IN2(~na26_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na347_1), .IN8(~na55_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x7y46     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6_1 ( .OUT(na6_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(na164_2), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a6_2 ( .OUT(na6_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a6_4 ( .OUT(na6_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(na164_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a6_5 ( .OUT(na6_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na6_2_i) );
// C_ORAND/D///      x11y38     80'h00_FE00_00_0000_0888_FEC3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1_i), .IN1(1'b0), .IN2(~na115_2), .IN3(1'b0), .IN4(na108_1), .IN5(na65_1), .IN6(na8_1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_2 ( .OUT(na8_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na8_1_i) );
// C_AND/D//AND/D      x22y37     80'h00_FE00_80_0000_0C88_4CAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9_1 ( .OUT(na9_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na315_2), .IN7(~na9_2), .IN8(na489_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a9_2 ( .OUT(na9_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na9_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9_4 ( .OUT(na9_2_i), .IN1(1'b1), .IN2(na115_2), .IN3(na386_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a9_5 ( .OUT(na9_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na9_2_i) );
// C_MX2b/D///      x16y45     80'h00_FE00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a10_1 ( .OUT(na10_1_i), .IN1(1'b1), .IN2(~na79_1), .IN3(1'b0), .IN4(1'b0), .IN5(na68_1), .IN6(na332_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a10_2 ( .OUT(na10_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na10_1_i) );
// C_MX4b/D///      x22y41     80'h00_FD00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a11_1 ( .OUT(na11_1_i), .IN1(na2_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na336_1), .IN5(1'b0), .IN6(1'b0), .IN7(na11_1), .IN8(na55_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a11_2 ( .OUT(na11_1), .CLK(~na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na11_1_i) );
// C_MX4b/D///      x13y36     80'h00_FD00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1_i), .IN1(na2_2), .IN2(1'b1), .IN3(1'b1), .IN4(na336_1), .IN5(na52_1), .IN6(na13_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a12_2 ( .OUT(na12_1), .CLK(~na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na12_1_i) );
// C_MX2a////      x15y40     80'h00_0018_00_0040_0C8C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1), .IN1(1'b0), .IN2(1'b0), .IN3(na59_1), .IN4(~na349_1), .IN5(1'b1), .IN6(na26_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP*/D//AND*/D      x15y33     80'h00_FE00_80_0000_0387_393A
C_ICOMP    #(.CPE_CFG (9'b1_0000_0000)) 
           _a14_1 ( .OUT(na14_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na14_2), .IN6(~na463_2), .IN7(1'b0), .IN8(na336_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a14_2 ( .OUT(na14_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na14_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a14_4 ( .OUT(na14_2_i), .IN1(na464_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na336_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a14_5 ( .OUT(na14_2), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na14_2_i) );
// C_AND/D///      x23y40     80'h00_FE00_00_0000_0888_2F22
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a15_1 ( .OUT(na15_1_i), .IN1(na103_1), .IN2(~na8_1), .IN3(na11_1), .IN4(~na60_1), .IN5(1'b1), .IN6(1'b1), .IN7(na58_2),
                    .IN8(~na61_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a15_2 ( .OUT(na15_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na15_1_i) );
// C_///AND/D      x7y44     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a18_4 ( .OUT(na18_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(1'b1), .IN4(na153_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a18_5 ( .OUT(na18_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na18_2_i) );
// C_AND/D//AND/D      x8y46     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a19_1 ( .OUT(na19_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(1'b1), .IN8(na162_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a19_2 ( .OUT(na19_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na19_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a19_4 ( .OUT(na19_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(1'b1), .IN4(na162_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a19_5 ( .OUT(na19_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na19_2_i) );
// C_AND/D//AND/D      x6y45     80'h00_FE00_80_0000_0C88_CC5C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a20_1 ( .OUT(na20_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(1'b1), .IN8(na153_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a20_2 ( .OUT(na20_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na20_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a20_4 ( .OUT(na20_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(~na20_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a20_5 ( .OUT(na20_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na20_2_i) );
// C_AND/D//AND/D      x7y42     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(na144_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a22_2 ( .OUT(na22_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na22_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a22_4 ( .OUT(na22_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(na144_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a22_5 ( .OUT(na22_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na22_2_i) );
// C_AND/D//AND/D      x22y45     80'h00_FE00_80_0000_0C88_ACCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a23_1 ( .OUT(na23_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na115_2), .IN7(na352_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a23_2 ( .OUT(na23_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na23_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a23_4 ( .OUT(na23_2_i), .IN1(1'b1), .IN2(na115_2), .IN3(1'b1), .IN4(na354_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a23_5 ( .OUT(na23_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na23_2_i) );
// C_AND/D///      x15y44     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a24_1 ( .OUT(na24_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na115_2), .IN7(na353_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a24_2 ( .OUT(na24_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na24_1_i) );
// C_AND/D//ORAND/D      x21y36     80'h00_FE00_80_0000_0C88_82EC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a26_1 ( .OUT(na26_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na493_2), .IN6(~na26_2), .IN7(na490_2), .IN8(na31_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a26_2 ( .OUT(na26_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na26_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a26_4 ( .OUT(na26_2_i), .IN1(1'b0), .IN2(na115_2), .IN3(na9_1), .IN4(na468_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a26_5 ( .OUT(na26_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na26_2_i) );
// C_AND/D//AND/D      x18y36     80'h00_FE00_80_0000_0C88_CCF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na115_2), .IN7(1'b1), .IN8(na355_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a27_2 ( .OUT(na27_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na27_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a27_4 ( .OUT(na27_2_i), .IN1(na351_1), .IN2(na115_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a27_5 ( .OUT(na27_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na27_2_i) );
// C_AND/D//AND/D      x21y44     80'h00_FE00_80_0000_0C88_F8CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a28_1 ( .OUT(na28_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na356_1), .IN6(na115_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a28_2 ( .OUT(na28_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na28_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a28_4 ( .OUT(na28_2_i), .IN1(1'b1), .IN2(na115_2), .IN3(1'b1), .IN4(na395_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a28_5 ( .OUT(na28_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na28_2_i) );
// C_///AND/D      x20y41     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a29_4 ( .OUT(na29_2_i), .IN1(1'b1), .IN2(na115_2), .IN3(na357_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a29_5 ( .OUT(na29_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na29_2_i) );
// C_AND/D//AND/D      x14y46     80'h00_FE00_80_0000_0C88_2AAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a30_1 ( .OUT(na30_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na126_1), .IN6(1'b1), .IN7(na110_1), .IN8(~na30_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a30_2 ( .OUT(na30_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na30_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a30_4 ( .OUT(na30_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na10_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a30_5 ( .OUT(na30_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na30_2_i) );
// C_ORAND/D//AND/D      x24y38     80'h00_FE00_80_0000_0C88_ECC4
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a31_1 ( .OUT(na31_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na115_2), .IN7(na472_2), .IN8(na31_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a31_2 ( .OUT(na31_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na31_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a31_4 ( .OUT(na31_2_i), .IN1(~na76_1), .IN2(na115_2), .IN3(1'b1), .IN4(na481_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a31_5 ( .OUT(na31_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na31_2_i) );
// C_AND/D//AND/D      x17y44     80'h00_FE00_80_0000_0C88_83CF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_1 ( .OUT(na33_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na33_2), .IN7(na39_2), .IN8(na51_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a33_2 ( .OUT(na33_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na33_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a33_4 ( .OUT(na33_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na51_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a33_5 ( .OUT(na33_2), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na33_2_i) );
// C_ORAND/D///      x17y41     80'h00_FE00_00_0000_0888_FE5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a35_1 ( .OUT(na35_1_i), .IN1(1'b0), .IN2(na488_2), .IN3(~na39_2), .IN4(1'b0), .IN5(na35_1), .IN6(na15_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a35_2 ( .OUT(na35_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na35_1_i) );
// C_AND/D///      x16y46     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na361_1), .IN7(1'b1), .IN8(na108_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a36_2 ( .OUT(na36_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na36_1_i) );
// C_///AND/      x13y39     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a37_4 ( .OUT(na37_2), .IN1(na80_1), .IN2(na8_1), .IN3(na58_2), .IN4(na74_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//ORAND/D      x24y41     80'h00_FE00_80_0000_0C88_AAEC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_1 ( .OUT(na39_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na130_2), .IN6(1'b1), .IN7(na39_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a39_2 ( .OUT(na39_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na39_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a39_4 ( .OUT(na39_2_i), .IN1(1'b0), .IN2(na488_2), .IN3(na39_2), .IN4(na363_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a39_5 ( .OUT(na39_2), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na39_2_i) );
// C_///AND/D      x19y42     80'h00_F600_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a40_4 ( .OUT(na40_2_i), .IN1(1'b1), .IN2(~na41_1), .IN3(1'b1), .IN4(na459_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a40_5 ( .OUT(na40_2), .CLK(na335_1), .EN(~na134_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na40_2_i) );
// C_ORAND////      x19y42     80'h00_0018_00_0000_0C88_A7FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a41_1 ( .OUT(na41_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na477_2), .IN6(~na50_1), .IN7(na39_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x12y45     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a42_1 ( .OUT(na42_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na113_1), .IN6(na492_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a42_2 ( .OUT(na42_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na42_1_i) );
// C_///AND/D      x22y48     80'h00_F600_80_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a43_4 ( .OUT(na43_2_i), .IN1(1'b1), .IN2(~na41_1), .IN3(na457_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a43_5 ( .OUT(na43_2), .CLK(na335_1), .EN(~na134_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na43_2_i) );
// C_AND/D///      x21y45     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a44_1 ( .OUT(na44_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na126_1), .IN6(1'b1), .IN7(1'b1), .IN8(na345_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a44_2 ( .OUT(na44_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na44_1_i) );
// C_AND/D///      x24y46     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na126_1), .IN6(na346_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a45_2 ( .OUT(na45_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na45_1_i) );
// C_///AND/D      x11y36     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a46_4 ( .OUT(na46_2_i), .IN1(na126_1), .IN2(na205_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a46_5 ( .OUT(na46_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na46_2_i) );
// C_AND/D///      x24y48     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a47_1 ( .OUT(na47_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na40_2), .IN7(na39_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a47_2 ( .OUT(na47_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na47_1_i) );
// C_///AND/D      x22y44     80'h00_FE00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a48_4 ( .OUT(na48_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na39_2), .IN4(na98_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a48_5 ( .OUT(na48_2), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na48_2_i) );
// C_///AND/D      x22y43     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a49_4 ( .OUT(na49_2_i), .IN1(1'b1), .IN2(na111_1), .IN3(na39_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a49_5 ( .OUT(na49_2), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na49_2_i) );
// C_ICOMP/D///      x27y46     80'h00_FE00_00_0000_0C88_A6FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a50_1 ( .OUT(na50_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na477_2), .IN6(~na50_1), .IN7(~na39_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a50_2 ( .OUT(na50_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na50_1_i) );
// C_///ORAND/D      x26y46     80'h00_FE00_80_0000_0C08_FFDC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a51_4 ( .OUT(na51_2_i), .IN1(1'b0), .IN2(na41_1), .IN3(~na58_2), .IN4(na51_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a51_5 ( .OUT(na51_2), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na51_2_i) );
// C_AND/D///      x17y37     80'h00_FD00_00_0000_0C88_1AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a52_1 ( .OUT(na52_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2_2), .IN6(1'b1), .IN7(~na336_1), .IN8(~na53_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a52_2 ( .OUT(na52_1), .CLK(~na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na52_1_i) );
// C_MX2b////      x22y40     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a53_1 ( .OUT(na53_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na468_2), .IN5(~na367_2), .IN6(1'b0), .IN7(~na59_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x15y45     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a54_1 ( .OUT(na54_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na126_1), .IN6(1'b1), .IN7(1'b1), .IN8(na30_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a54_2 ( .OUT(na54_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na54_1_i) );
// C_AND/D//AND/D      x20y36     80'h00_FE00_80_0000_0C88_C32F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na336_1), .IN7(1'b1), .IN8(na55_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a55_2 ( .OUT(na55_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na55_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a55_4 ( .OUT(na55_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na59_1), .IN4(~na336_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a55_5 ( .OUT(na55_2), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na55_2_i) );
// C_AND/D///      x14y42     80'h00_FE00_00_0000_0888_234A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a57_1 ( .OUT(na57_1_i), .IN1(na103_1), .IN2(1'b1), .IN3(~na11_1), .IN4(na61_1), .IN5(1'b1), .IN6(~na8_1), .IN7(na58_2),
                    .IN8(~na60_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a57_2 ( .OUT(na57_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na57_1_i) );
// C_///AND/D      x22y39     80'h00_FD00_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a58_4 ( .OUT(na58_2_i), .IN1(na2_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na336_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a58_5 ( .OUT(na58_2), .CLK(~na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na58_2_i) );
// C_AND/D//AND/D      x20y39     80'h00_FE00_80_0000_0C88_2F3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a59_1 ( .OUT(na59_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na59_2), .IN8(~na336_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a59_2 ( .OUT(na59_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na59_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a59_4 ( .OUT(na59_2_i), .IN1(1'b1), .IN2(na334_1), .IN3(1'b1), .IN4(~na336_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a59_5 ( .OUT(na59_2), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na59_2_i) );
// C_MX4b/D///      x12y40     80'h00_FD00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a60_1 ( .OUT(na60_1_i), .IN1(~na2_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na336_1), .IN5(1'b0), .IN6(1'b0), .IN7(na59_2), .IN8(na60_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a60_2 ( .OUT(na60_1), .CLK(~na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na60_1_i) );
// C_MX4b/D///      x16y38     80'h00_FD00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a61_1 ( .OUT(na61_1_i), .IN1(~na2_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na336_1), .IN5(1'b0), .IN6(1'b0), .IN7(na59_1), .IN8(na61_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a61_2 ( .OUT(na61_1), .CLK(~na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na61_1_i) );
// C_AND/D//AND/D      x24y43     80'h00_FE00_80_0000_0C88_F8AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a62_1 ( .OUT(na62_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na368_1), .IN6(na115_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a62_2 ( .OUT(na62_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na62_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a62_4 ( .OUT(na62_2_i), .IN1(1'b1), .IN2(na115_2), .IN3(na369_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a62_5 ( .OUT(na62_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na62_2_i) );
// C_AND/D//AND/D      x14y47     80'h00_FE00_80_0000_0C88_4AAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a64_1 ( .OUT(na64_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na126_1), .IN6(1'b1), .IN7(~na110_1), .IN8(na30_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a64_2 ( .OUT(na64_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na64_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a64_4 ( .OUT(na64_2_i), .IN1(na126_1), .IN2(1'b1), .IN3(na64_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a64_5 ( .OUT(na64_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na64_2_i) );
// C_AND/D///      x21y37     80'h00_FE00_00_0000_0888_8325
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a65_1 ( .OUT(na65_1_i), .IN1(~na103_1), .IN2(1'b1), .IN3(na58_2), .IN4(~na61_1), .IN5(1'b1), .IN6(~na8_1), .IN7(na11_1),
                    .IN8(na60_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a65_2 ( .OUT(na65_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na65_1_i) );
// C_AND/D//AND/D      x7y45     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_1 ( .OUT(na67_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(na157_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a67_2 ( .OUT(na67_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na67_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a67_4 ( .OUT(na67_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(na157_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a67_5 ( .OUT(na67_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na67_2_i) );
// C_AND/D///      x15y47     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a68_1 ( .OUT(na68_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na333_1), .IN6(na492_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a68_2 ( .OUT(na68_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na68_1_i) );
// C_///AND/D      x12y43     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a72_4 ( .OUT(na72_2_i), .IN1(1'b1), .IN2(na370_1), .IN3(1'b1), .IN4(na108_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a72_5 ( .OUT(na72_2), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na72_2_i) );
// C_AND////      x19y44     80'h00_0018_00_0000_0C88_28FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a73_1 ( .OUT(na73_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na80_1), .IN6(na8_1), .IN7(na58_2), .IN8(~na74_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a/D///      x14y48     80'h00_FE00_00_0040_0C0C_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a74_1 ( .OUT(na74_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na371_2), .IN4(na74_1), .IN5(1'b1), .IN6(~na8_1), .IN7(1'b1), .IN8(na108_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a74_2 ( .OUT(na74_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na74_1_i) );
// C_AND/D///      x13y43     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na372_1), .IN7(1'b1), .IN8(na108_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a75_2 ( .OUT(na75_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na75_1_i) );
// C_AND/D//AND/D      x17y39     80'h00_FE00_80_0000_0C88_CCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a76_1 ( .OUT(na76_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na115_2), .IN7(1'b1), .IN8(na373_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a76_2 ( .OUT(na76_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na76_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a76_4 ( .OUT(na76_2_i), .IN1(na76_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a76_5 ( .OUT(na76_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na76_2_i) );
// C_AND/D//AND/D      x19y48     80'h00_FE00_80_0000_0C88_ACF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a77_1 ( .OUT(na77_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na115_2), .IN7(na374_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a77_2 ( .OUT(na77_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na77_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a77_4 ( .OUT(na77_2_i), .IN1(na359_1), .IN2(na115_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a77_5 ( .OUT(na77_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na77_2_i) );
// C_AND/D//AND/D      x10y46     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(1'b1), .IN8(na155_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a78_2 ( .OUT(na78_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a78_4 ( .OUT(na78_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(1'b1), .IN4(na155_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a78_5 ( .OUT(na78_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_2_i) );
// C_AND/D///      x13y44     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a79_1 ( .OUT(na79_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na375_1), .IN7(1'b1), .IN8(na108_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a79_2 ( .OUT(na79_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na79_1_i) );
// C_ICOMP/D///      x21y41     80'h00_FE00_00_0000_0C88_C6FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na80_1), .IN6(~na81_2), .IN7(1'b0), .IN8(~na108_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a80_2 ( .OUT(na80_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na80_1_i) );
// C_///AND/      x19y44     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a81_4 ( .OUT(na81_2), .IN1(1'b1), .IN2(na8_1), .IN3(na58_2), .IN4(na74_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x10y45     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a84_1 ( .OUT(na84_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(na152_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a84_2 ( .OUT(na84_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na84_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a84_4 ( .OUT(na84_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(na152_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a84_5 ( .OUT(na84_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na84_2_i) );
// C_AND/D//AND/D      x7y43     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a87_1 ( .OUT(na87_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(1'b1), .IN8(na150_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a87_2 ( .OUT(na87_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na87_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a87_4 ( .OUT(na87_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(1'b1), .IN4(na150_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a87_5 ( .OUT(na87_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na87_2_i) );
// C_AND/D//AND/D      x10y43     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(na148_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a89_2 ( .OUT(na89_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a89_4 ( .OUT(na89_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(na148_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a89_5 ( .OUT(na89_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_2_i) );
// C_AND/D//AND/D      x13y41     80'h00_FE00_80_0000_0C88_CCF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na379_1), .IN7(1'b1), .IN8(na489_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a90_2 ( .OUT(na90_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na90_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a90_4 ( .OUT(na90_2_i), .IN1(na377_1), .IN2(na115_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a90_5 ( .OUT(na90_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na90_2_i) );
// C_///ICOMP/D      x21y40     80'h00_FE00_80_0000_0C08_FF9C
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a91_4 ( .OUT(na91_2_i), .IN1(1'b0), .IN2(~na115_2), .IN3(~na484_2), .IN4(~na468_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a91_5 ( .OUT(na91_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na91_2_i) );
// C_OR/D///      x19y35     80'h00_FE00_00_0000_0CEE_0B00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a92_1 ( .OUT(na92_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na381_1), .IN6(~na115_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a92_2 ( .OUT(na92_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na92_1_i) );
// C_///AND/D      x22y36     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a93_4 ( .OUT(na93_2_i), .IN1(1'b1), .IN2(na115_2), .IN3(na382_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a93_5 ( .OUT(na93_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na93_2_i) );
// C_AND/D///      x19y36     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a94_1 ( .OUT(na94_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na115_2), .IN7(1'b1), .IN8(na383_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a94_2 ( .OUT(na94_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na94_1_i) );
// C_AND/D//AND/D      x17y47     80'h00_FE00_80_0000_0C88_F8AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a96_1 ( .OUT(na96_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na384_1), .IN6(na115_2), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a96_2 ( .OUT(na96_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na96_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a96_4 ( .OUT(na96_2_i), .IN1(1'b1), .IN2(na115_2), .IN3(na391_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a96_5 ( .OUT(na96_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na96_2_i) );
// C_///AND/D      x22y46     80'h00_F600_80_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a98_4 ( .OUT(na98_2_i), .IN1(1'b1), .IN2(~na41_1), .IN3(na460_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a98_5 ( .OUT(na98_2), .CLK(na335_1), .EN(~na134_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na98_2_i) );
// C_ICOMP/D///      x20y35     80'h00_FE00_00_0000_0C88_6CFF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a100_1 ( .OUT(na100_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na115_2), .IN7(na100_1), .IN8(~na467_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a100_2 ( .OUT(na100_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na100_1_i) );
// C_AND/D//AND/D      x20y34     80'h00_FE00_80_0000_0C88_F8CC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a102_1 ( .OUT(na102_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na389_1), .IN6(na115_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a102_2 ( .OUT(na102_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na102_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a102_4 ( .OUT(na102_2_i), .IN1(1'b1), .IN2(na115_2), .IN3(1'b1), .IN4(na388_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a102_5 ( .OUT(na102_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na102_2_i) );
// C_MX4b/D///      x13y37     80'h00_FD00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_1 ( .OUT(na103_1_i), .IN1(na2_2), .IN2(1'b1), .IN3(1'b1), .IN4(na336_1), .IN5(na103_1), .IN6(na476_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a103_2 ( .OUT(na103_1), .CLK(~na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na103_1_i) );
// C_AND/D//AND/D      x6y46     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a106_1 ( .OUT(na106_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(1'b1), .IN8(na146_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a106_2 ( .OUT(na106_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na106_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a106_4 ( .OUT(na106_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(1'b1), .IN4(na146_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a106_5 ( .OUT(na106_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na106_2_i) );
// C_ORAND/D///      x18y44     80'h00_FE00_00_0000_0888_EF3C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a108_1 ( .OUT(na108_1_i), .IN1(1'b0), .IN2(na350_2), .IN3(1'b0), .IN4(~na57_1), .IN5(1'b1), .IN6(1'b1), .IN7(na247_2), .IN8(na108_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a108_2 ( .OUT(na108_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na108_1_i) );
// C_MX2b/D///      x16y47     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a110_1 ( .OUT(na110_1_i), .IN1(na126_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na10_1), .IN8(na30_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a110_2 ( .OUT(na110_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na110_1_i) );
// C_MX2b/D///      x23y44     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a111_1 ( .OUT(na111_1_i), .IN1(1'b1), .IN2(na41_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na461_1), .IN8(na43_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a111_2 ( .OUT(na111_1), .CLK(na335_1), .EN(~na134_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na111_1_i) );
// C_AND/D//AND/D      x6y47     80'h00_FE00_80_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a112_1 ( .OUT(na112_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(1'b1), .IN8(na166_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a112_2 ( .OUT(na112_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na112_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a112_4 ( .OUT(na112_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(1'b1), .IN4(na166_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a112_5 ( .OUT(na112_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na112_2_i) );
// C_AND/D//AND/D      x9y45     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a113_1 ( .OUT(na113_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na350_2), .IN7(na160_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a113_2 ( .OUT(na113_1), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na113_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a113_4 ( .OUT(na113_2_i), .IN1(1'b1), .IN2(na350_2), .IN3(na160_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a113_5 ( .OUT(na113_2), .CLK(na205_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na113_2_i) );
// C_///ORAND/D      x19y38     80'h00_FE00_80_0000_0C08_FFCE
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a115_4 ( .OUT(na115_2_i), .IN1(na37_2), .IN2(na115_2), .IN3(1'b0), .IN4(na108_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a115_5 ( .OUT(na115_2), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na115_2_i) );
// C_MX2b/D///      x18y47     80'h00_F600_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a116_1 ( .OUT(na116_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na23_2), .IN8(~na491_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a116_2 ( .OUT(na116_1), .CLK(na335_1), .EN(~na133_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na116_1_i) );
// C_MX2b/D///      x17y46     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a117_1 ( .OUT(na117_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na177_1), .IN8(na494_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a117_2 ( .OUT(na117_1), .CLK(na335_1), .EN(~na133_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na117_1_i) );
// C_MX2b/D///      x18y46     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a118_1 ( .OUT(na118_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na177_2), .IN8(na495_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a118_2 ( .OUT(na118_1), .CLK(na335_1), .EN(~na133_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na118_1_i) );
// C_MX2b/D///      x20y45     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a119_1 ( .OUT(na119_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na498_2), .IN8(na170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a119_2 ( .OUT(na119_1), .CLK(na335_1), .EN(~na133_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na119_1_i) );
// C_MX2b/D///      x19y46     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a120_1 ( .OUT(na120_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na499_2), .IN8(na170_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a120_2 ( .OUT(na120_1), .CLK(na335_1), .EN(~na133_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na120_1_i) );
// C_MX2b/D///      x20y46     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a121_1 ( .OUT(na121_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na181_1), .IN8(na496_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a121_2 ( .OUT(na121_1), .CLK(na335_1), .EN(~na133_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na121_1_i) );
// C_MX2b/D///      x21y47     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a122_1 ( .OUT(na122_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na181_2), .IN8(na497_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a122_2 ( .OUT(na122_1), .CLK(na335_1), .EN(~na133_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na122_1_i) );
// C_MX2b/D///      x22y47     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a123_1 ( .OUT(na123_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na500_2), .IN8(na174_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a123_2 ( .OUT(na123_1), .CLK(na335_1), .EN(~na133_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na123_1_i) );
// C_MX2b/D///      x21y42     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a124_1 ( .OUT(na124_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na501_2), .IN8(na174_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a124_2 ( .OUT(na124_1), .CLK(na335_1), .EN(~na133_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na124_1_i) );
// C_AND/D///      x18y43     80'h00_FE00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a125_1 ( .OUT(na125_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na393_1), .IN8(na108_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a125_2 ( .OUT(na125_1), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na125_1_i) );
// C_ORAND/D///      x11y45     80'h00_FE00_00_0000_0888_FE3C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a126_1 ( .OUT(na126_1_i), .IN1(1'b0), .IN2(na350_2), .IN3(1'b0), .IN4(~na57_1), .IN5(na126_1), .IN6(na248_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a126_2 ( .OUT(na126_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na126_1_i) );
// C_///AND/D      x21y43     80'h00_F600_80_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a130_4 ( .OUT(na130_2_i), .IN1(1'b1), .IN2(~na41_1), .IN3(1'b1), .IN4(na458_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a130_5 ( .OUT(na130_2), .CLK(na335_1), .EN(~na134_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na130_2_i) );
// C_AND/D//AND/D      x22y35     80'h00_FE00_80_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a131_1 ( .OUT(na131_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na115_2), .IN7(na396_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a131_2 ( .OUT(na131_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na131_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a131_4 ( .OUT(na131_2_i), .IN1(1'b1), .IN2(na115_2), .IN3(na378_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a131_5 ( .OUT(na131_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na131_2_i) );
// C_ORAND////      x23y45     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a133_1 ( .OUT(na133_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na475_2), .IN6(~na26_2), .IN7(1'b0), .IN8(~na473_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x22y46     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a134_1 ( .OUT(na134_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na41_1), .IN7(~na58_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x13y45     80'h00_0018_00_0040_0C05_2000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(na54_1), .IN2(1'b0), .IN3(na64_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na125_1), .IN8(~na36_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x18y48     80'h00_FE00_80_0000_0C08_FFEA
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a139_4 ( .OUT(na139_2_i), .IN1(na126_1), .IN2(1'b0), .IN3(na401_2), .IN4(na139_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a139_5 ( .OUT(na139_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na139_2_i) );
// C_MX2b////      x22y38     80'h00_0018_00_0040_0AC8_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a140_1 ( .OUT(na140_1), .IN1(1'b1), .IN2(~na26_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na402_1), .IN8(~na55_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x18y30     80'h00_FD00_00_0000_0888_3F7E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a141_1 ( .OUT(na141_1_i), .IN1(na2_2), .IN2(na1_1), .IN3(~na462_2), .IN4(~na140_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0), .IN8(~na336_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a141_2 ( .OUT(na141_1), .CLK(~na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na141_1_i) );
// C_ADDF2///ADDF2/      x8y39     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a144_1 ( .OUT(na144_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na22_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na166_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a144_4 ( .OUT(na144_2), .COUTY1(na144_4), .IN1(1'b1), .IN2(na22_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na22_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na166_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x8y40     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a146_1 ( .OUT(na146_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na106_2),
                     .CINX(1'b0), .CINY1(na144_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a146_4 ( .OUT(na146_2), .COUTY1(na146_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na106_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na106_2), .CINX(1'b0), .CINY1(na144_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x8y41     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a148_1 ( .OUT(na148_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na89_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na146_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a148_4 ( .OUT(na148_2), .COUTY1(na148_4), .IN1(1'b0), .IN2(1'b0), .IN3(na89_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na89_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na146_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x8y42     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a150_1 ( .OUT(na150_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na87_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na148_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a150_4 ( .OUT(na150_2), .COUTY1(na150_4), .IN1(na87_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na87_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na148_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x8y43     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a152_1 ( .OUT(na152_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na84_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na150_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a152_4 ( .OUT(na152_2), .COUTY1(na152_4), .IN1(1'b0), .IN2(1'b0), .IN3(na84_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na84_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na150_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x8y34     80'h00_0078_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a153_1 ( .OUT(na153_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na18_2), .IN7(na20_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na167_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a153_4 ( .OUT(na153_2), .COUTY1(na153_4), .IN1(1'b0), .IN2(1'b0), .IN3(na20_1), .IN4(1'b1), .IN5(1'b1), .IN6(na18_2), .IN7(na20_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na167_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x8y44     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a155_1 ( .OUT(na155_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na78_2),
                     .CINX(1'b0), .CINY1(na152_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a155_4 ( .OUT(na155_2), .COUTY1(na155_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na78_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na78_2), .CINX(1'b0), .CINY1(na152_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x8y45     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a157_1 ( .OUT(na157_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na67_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na155_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a157_4 ( .OUT(na157_2), .IN1(na67_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na67_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na155_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x8y35     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a160_1 ( .OUT(na160_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na113_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na153_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a160_4 ( .OUT(na160_2), .COUTY1(na160_4), .IN1(na113_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na113_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na153_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x8y36     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a162_1 ( .OUT(na162_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na19_2),
                     .CINX(1'b0), .CINY1(na160_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a162_4 ( .OUT(na162_2), .COUTY1(na162_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na19_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na19_2), .CINX(1'b0), .CINY1(na160_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x8y37     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a164_1 ( .OUT(na164_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na6_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na162_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a164_4 ( .OUT(na164_2), .COUTY1(na164_4), .IN1(1'b1), .IN2(na6_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na6_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na162_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x8y38     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a166_1 ( .OUT(na166_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na112_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na164_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a166_4 ( .OUT(na166_2), .COUTY1(na166_4), .IN1(1'b0), .IN2(1'b0), .IN3(na112_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na112_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na164_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x8y33     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a167_2 ( .OUT(na167_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a167_6 ( .COUTY1(na167_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na167_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x18y39     80'h00_0078_00_0020_0C66_ACC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a168_1 ( .OUT(na168_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na117_1), .IN7(na116_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na176_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a168_4 ( .OUT(na168_2), .COUTY1(na168_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na118_1), .IN5(1'b1), .IN6(na117_1), .IN7(na116_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na176_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x18y40     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a170_1 ( .OUT(na170_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na119_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na168_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a170_4 ( .OUT(na170_2), .COUTY1(na170_4), .IN1(1'b1), .IN2(na120_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na119_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na168_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x18y41     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a172_1 ( .OUT(na172_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na121_1),
                     .CINX(1'b0), .CINY1(na170_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a172_4 ( .OUT(na172_2), .COUTY1(na172_4), .IN1(na122_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na121_1), .CINX(1'b0), .CINY1(na170_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x18y42     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a174_1 ( .OUT(na174_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na123_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na172_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a174_4 ( .OUT(na174_2), .IN1(1'b1), .IN2(na124_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na123_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na172_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x18y38     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a176_2 ( .OUT(na176_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a176_6 ( .COUTY1(na176_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na176_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x16y41     80'h00_0078_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a177_1 ( .OUT(na177_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na24_1), .IN7(na23_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na185_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a177_4 ( .OUT(na177_2), .COUTY1(na177_4), .IN1(1'b0), .IN2(1'b0), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(na24_1), .IN7(na23_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na185_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x16y42     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a179_1 ( .OUT(na179_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na28_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na177_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a179_4 ( .OUT(na179_2), .COUTY1(na179_4), .IN1(1'b1), .IN2(na28_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na28_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na177_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x16y43     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a181_1 ( .OUT(na181_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na96_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na179_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a181_4 ( .OUT(na181_2), .COUTY1(na181_4), .IN1(na96_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na96_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na179_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x16y44     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a183_1 ( .OUT(na183_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na77_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na181_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a183_4 ( .OUT(na183_2), .IN1(1'b1), .IN2(na77_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na77_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na181_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x16y40     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a185_2 ( .OUT(na185_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a185_6 ( .COUTY1(na185_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na185_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x15y36     80'h00_0078_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a186_1 ( .OUT(na186_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na91_2), .IN7(na62_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na194_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a186_4 ( .OUT(na186_2), .COUTY1(na186_4), .IN1(1'b0), .IN2(1'b0), .IN3(na62_1), .IN4(1'b1), .IN5(1'b1), .IN6(na91_2), .IN7(na62_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na194_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x15y37     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a188_1 ( .OUT(na188_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na27_2),
                     .CINX(1'b0), .CINY1(na186_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a188_4 ( .OUT(na188_2), .COUTY1(na188_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na27_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na27_2), .CINX(1'b0), .CINY1(na186_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x15y38     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a190_1 ( .OUT(na190_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na76_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na188_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a190_4 ( .OUT(na190_2), .COUTY1(na190_4), .IN1(1'b0), .IN2(1'b0), .IN3(na29_2), .IN4(1'b1), .IN5(na76_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na188_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x15y39     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a192_1 ( .OUT(na192_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na90_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na190_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a192_4 ( .OUT(na192_2), .IN1(na90_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na90_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na190_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x15y35     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a194_2 ( .OUT(na194_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a194_6 ( .COUTY1(na194_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na194_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x20y29     80'h00_0078_00_0020_0C66_CAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a195_1 ( .OUT(na195_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na487_2), .IN6(1'b1), .IN7(1'b1), .IN8(na102_2),
                     .CINX(1'b0), .CINY1(na344_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a195_4 ( .OUT(na195_2), .COUTY1(na195_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na102_1), .IN5(na487_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na102_2), .CINX(1'b0), .CINY1(na344_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x20y30     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a197_1 ( .OUT(na197_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na131_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na195_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a197_4 ( .OUT(na197_2), .COUTY1(na197_4), .IN1(1'b0), .IN2(1'b0), .IN3(na131_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na131_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na195_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x20y31     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a199_1 ( .OUT(na199_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na93_2),
                     .CINX(1'b0), .CINY1(na197_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a199_4 ( .OUT(na199_2), .COUTY1(na199_4), .IN1(na92_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na93_2), .CINX(1'b0), .CINY1(na197_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x20y32     80'h00_0078_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a201_1 ( .OUT(na201_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na94_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na199_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a201_4 ( .OUT(na201_2), .IN1(1'b0), .IN2(1'b0), .IN3(na9_2), .IN4(1'b1), .IN5(1'b1), .IN6(na94_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na199_4), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0014_0016)) 
           _a205 ( .GLB0(na205_1), .GLB1(na205_2), .GLB2(_d0), .GLB3(_d1), .CLK_FB0(_d2), .CLK_FB1(_d3), .CLK_FB2(_d4), .CLK_FB3(_d5),
                   .CLK0_0(na340_6), .CLK0_90(na340_5), .CLK0_180(na340_4), .CLK0_270(na340_3), .CLK0_BYP(1'b0), .CLK1_0(na339_6),
                   .CLK1_90(na339_5), .CLK1_180(na339_4), .CLK1_270(na339_3), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0),
                   .CLK2_270(1'b0), .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0),
                   .USR_GLB0(1'b0), .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0),
                   .USR_FB3(1'b0) );
// C_///AND/D      x14y43     80'h00_FE00_80_0000_0C08_FF3F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a247_4 ( .OUT(na247_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na108_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a247_5 ( .OUT(na247_2), .CLK(na335_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na247_2_i) );
// C_AND/D///      x15y48     80'h00_FE00_00_0000_0C88_F5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a248_1 ( .OUT(na248_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na126_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a248_2 ( .OUT(na248_1), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na248_1_i) );
// C_///AND/D      x19y36     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a315_4 ( .OUT(na315_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na9_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a315_5 ( .OUT(na315_2), .CLK(na205_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na315_2_i) );
// C_MX4b////      x17y48     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a332_1 ( .OUT(na332_1), .IN1(na75_1), .IN2(1'b1), .IN3(~na72_2), .IN4(1'b1), .IN5(na44_1), .IN6(na46_2), .IN7(na42_1), .IN8(na45_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a333 ( .Y(na333_1), .I(clk) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a334 ( .Y(na334_1), .I(i_mosi_ILA) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a335 ( .Y(na335_1), .I(i_sclk_ILA) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a336 ( .Y(na336_1), .I(i_ss_ILA) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a337 ( .O(led), .A(na403_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a338 ( .O(o_miso_ILA), .A(na404_10) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_0C_08_0C_20_82)) 
           _a339 ( .USR_PLL_LOCKED_STDY(_d6), .USR_PLL_LOCKED(_d7), .CLK270(na339_3), .CLK180(na339_4), .CLK90(na339_5), .CLK0(na339_6),
                   .CLK_REF_OUT(_d8), .CLK_REF(na348_2), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_50_08_0C_20_82)) 
           _a340 ( .USR_PLL_LOCKED_STDY(_d9), .USR_PLL_LOCKED(_d10), .CLK270(na340_3), .CLK180(na340_4), .CLK90(na340_5), .CLK0(na340_6),
                   .CLK_REF_OUT(_d11), .CLK_REF(na348_1), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_08_20_0A_03_00_00_61_03_13_00_00_00_00_00_13_23_00_00_23_00_00),
             .INIT_00(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_01(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_02(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_03(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_04(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_05(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a341 ( .DOA({_d12, _d13, _d14, _d15, _d16, _d17, _d18, _d19, _d20, _d21, _d22, _d23, _d24, _d25, _d26, _d27, _d28, _d29,
                  _d30, _d31, _d32, _d33, _d34, _d35, _d36, _d37, _d38, _d39, _d40, _d41, _d42, _d43, _d44, _d45, _d46, _d47, _d48,
                  _d49, _d50, _d51}),
                   .DOAX({_d52, _d53, _d54, _d55, _d56, _d57, _d58, _d59, _d60, _d61, _d62, _d63, _d64, _d65, _d66, _d67, _d68, _d69,
                  _d70, _d71, _d72, _d73, _d74, _d75, _d76, _d77, _d78, _d79, _d80, _d81, _d82, _d83, _d84, _d85, _d86, _d87, _d88,
                  _d89, _d90, _d91}),
                   .DOB({_d92, _d93, _d94, _d95, _d96, _d97, _d98, _d99, _d100, _d101, _d102, _d103, _d104, _d105, _d106, na341_96,
                  na341_97, na341_98, na341_99, na341_100, _d107, _d108, _d109, _d110, _d111, _d112, _d113, _d114, _d115, _d116, _d117,
                  _d118, _d119, _d120, _d121, _d122, _d123, _d124, _d125, _d126}),
                   .DOBX({_d127, _d128, _d129, _d130, _d131, _d132, _d133, _d134, _d135, _d136, _d137, _d138, _d139, _d140, _d141,
                  _d142, _d143, _d144, _d145, _d146, _d147, _d148, _d149, _d150, _d151, _d152, _d153, _d154, _d155, _d156, _d157, _d158,
                  _d159, _d160, _d161, _d162, _d163, _d164, _d165, _d166}),
                   .ECC1B_ERRA({_d167, _d168, _d169, _d170}),
                   .ECC1B_ERRB({_d171, _d172, _d173, _d174}),
                   .ECC2B_ERRA({_d175, _d176, _d177, _d178}),
                   .ECC2B_ERRB({_d179, _d180, _d181, _d182}),
                   .FORW_CAS_WRAO(_d183), .FORW_CAS_WRBO(_d184), .FORW_CAS_BMAO(_d185), .FORW_CAS_BMBO(_d186), .FORW_CAS_RDAO(_d187),
                   .FORW_CAS_RDBO(_d188), .FORW_UADDRAO({_d189, _d190, _d191, _d192, _d193, _d194, _d195, _d196, _d197, _d198, _d199,
                  _d200, _d201, _d202, _d203, _d204}),
                   .FORW_LADDRAO({_d205, _d206, _d207, _d208, _d209, _d210, _d211, _d212, _d213, _d214, _d215, _d216, _d217, _d218,
                  _d219, _d220}),
                   .FORW_UADDRBO({_d221, _d222, _d223, _d224, _d225, _d226, _d227, _d228, _d229, _d230, _d231, _d232, _d233, _d234,
                  _d235, _d236}),
                   .FORW_LADDRBO({_d237, _d238, _d239, _d240, _d241, _d242, _d243, _d244, _d245, _d246, _d247, _d248, _d249, _d250,
                  _d251, _d252}),
                   .FORW_UA0CLKO(_d253), .FORW_UA0ENO(_d254), .FORW_UA0WEO(_d255), .FORW_LA0CLKO(_d256), .FORW_LA0ENO(_d257), .FORW_LA0WEO(_d258),
                   .FORW_UA1CLKO(_d259), .FORW_UA1ENO(_d260), .FORW_UA1WEO(_d261), .FORW_LA1CLKO(_d262), .FORW_LA1ENO(_d263), .FORW_LA1WEO(_d264),
                   .FORW_UB0CLKO(_d265), .FORW_UB0ENO(_d266), .FORW_UB0WEO(_d267), .FORW_LB0CLKO(_d268), .FORW_LB0ENO(_d269), .FORW_LB0WEO(_d270),
                   .FORW_UB1CLKO(_d271), .FORW_UB1ENO(_d272), .FORW_UB1WEO(_d273), .FORW_LB1CLKO(_d274), .FORW_LB1ENO(_d275), .FORW_LB1WEO(_d276),
                   .CLOCKA({_d277, _d278, _d279, _d280}),
                   .CLOCKB({_d281, _d282, _d283, _d284}),
                   .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .CLKB({1'b1, na358_9, 1'b1, 1'b1}),
                   .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .GLWEA({1'b1, na360_10, 1'b1, 1'b1}),
                   .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA1({na362_10, na364_9, na365_10, na366_9, na376_10, na380_9, na385_10, na387_9, na390_10, na392_9, na394_10,
                  na397_9, na398_10, na399_9, na400_10, na405_9}),
                   .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .ADDRB1({na406_10, na407_9, na408_10, na409_9, na410_10, na411_9, na412_10, na413_9, na414_10, na415_9, na416_10,
                  na417_9, na418_10, na419_9, na420_10, na421_9}),
                   .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .DIA({na422_10, na423_9, na424_10, na425_9, na426_10, na427_9, na428_10, na429_9, na430_10, na431_9, na432_10, na433_9,
                  na434_10, na435_9, na436_10, na437_9, na438_10, na439_9, na440_10, na441_9, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .WEA({na442_10, na443_9, na444_10, na445_9, na446_10, na447_9, na448_10, na449_9, na450_10, na451_9, na452_10, na453_9,
                  na454_10, na455_9, na456_10, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1}),
                   .CLOCK1(na205_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                   .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                  1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                   .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                   .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                   .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                   .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
CC_USR_RSTN            _a342 ( .USR_RSTN(na342_1) );
// C_///OR/      x18y38     80'h00_0060_00_0000_0C0E_FF3D
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a343_4 ( .OUT(na343_2), .IN1(~na2_2), .IN2(na4_1), .IN3(1'b0), .IN4(~na5_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x20y28     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a344_2 ( .OUT(na344_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a344_6 ( .COUTY1(na344_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na344_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x46y128     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a345_2 ( .OUT(na345_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na339_3), .CP_O(1'b0) );
// C_/RAM_I1///      x45y128     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a346_2 ( .OUT(na346_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na339_4), .CP_O(1'b0) );
// C_AND////      x24y45     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a347_1 ( .OUT(na347_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na35_1), .IN6(1'b1), .IN7(~na39_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a348 ( .PCLK0(na348_1), .PCLK1(na348_2), .PCLK2(_d285), .PCLK3(_d286), .CLK0(na333_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0),
                   .SER_CLK(1'b0), .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_AND////      x24y40     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a349_1 ( .OUT(na349_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na39_2), .IN8(~na48_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x1y66     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a350_5 ( .OUT(na350_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na342_1), .CP_O(1'b0) );
// C_MX2b////      x23y39     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a351_1 ( .OUT(na351_1), .IN1(1'b1), .IN2(na26_2), .IN3(1'b0), .IN4(1'b0), .IN5(na188_1), .IN6(na470_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x14y45     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a352_1 ( .OUT(na352_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na468_2), .IN5(na466_2), .IN6(1'b0), .IN7(na62_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x20y37     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a353_1 ( .OUT(na353_1), .IN1(1'b1), .IN2(na26_2), .IN3(1'b0), .IN4(1'b0), .IN5(na479_2), .IN6(na24_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x20y38     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a354_1 ( .OUT(na354_1), .IN1(1'b1), .IN2(~na26_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na23_2), .IN8(na485_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x14y36     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a355_1 ( .OUT(na355_1), .IN1(1'b1), .IN2(na26_2), .IN3(1'b0), .IN4(1'b0), .IN5(na188_2), .IN6(na469_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x19y45     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a356_1 ( .OUT(na356_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na468_2), .IN5(1'b0), .IN6(na28_1), .IN7(1'b0), .IN8(na27_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x14y37     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a357_1 ( .OUT(na357_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na468_2), .IN5(1'b0), .IN6(na190_2), .IN7(1'b0), .IN8(na471_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y57     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a358_1 ( .OUT(na358_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na335_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a358_6 ( .RAM_O1(na358_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na358_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x17y43     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a359_1 ( .OUT(na359_1), .IN1(1'b1), .IN2(na26_2), .IN3(1'b0), .IN4(1'b0), .IN5(na90_2), .IN6(na77_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x27y57     80'h08_0060_00_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a360_4 ( .OUT(na360_2), .IN1(1'b1), .IN2(~na26_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a360_6 ( .RAM_O2(na360_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na360_2), .COMP_OUT(1'b0) );
// C_MX2b////      x17y50     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a361_1 ( .OUT(na361_1), .IN1(na37_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na474_2), .IN8(na61_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a362_4 ( .OUT(na362_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a362_6 ( .RAM_O2(na362_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na362_2), .COMP_OUT(1'b0) );
// C_///AND/      x20y40     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a363_4 ( .OUT(na363_2), .IN1(na35_1), .IN2(1'b1), .IN3(na58_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a364_1 ( .OUT(na364_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a364_6 ( .RAM_O1(na364_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na364_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a365_4 ( .OUT(na365_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a365_6 ( .RAM_O2(na365_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na365_2), .COMP_OUT(1'b0) );
// C_AND////      x28y63     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a366_1 ( .OUT(na366_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na77_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a366_6 ( .RAM_O1(na366_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na366_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x19y39     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a367_4 ( .OUT(na367_2), .IN1(na475_2), .IN2(1'b1), .IN3(na49_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x13y35     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a368_1 ( .OUT(na368_1), .IN1(1'b1), .IN2(~na26_2), .IN3(1'b0), .IN4(1'b0), .IN5(na478_2), .IN6(na186_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x16y37     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a369_1 ( .OUT(na369_1), .IN1(1'b1), .IN2(~na26_2), .IN3(1'b0), .IN4(1'b0), .IN5(na479_2), .IN6(na186_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x13y48     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a370_1 ( .OUT(na370_1), .IN1(1'b1), .IN2(na73_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na72_2), .IN8(na60_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x18y45     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a371_4 ( .OUT(na371_2), .IN1(1'b0), .IN2(1'b0), .IN3(na58_2), .IN4(na74_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x15y46     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a372_1 ( .OUT(na372_1), .IN1(1'b1), .IN2(na73_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na480_2), .IN8(na61_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x14y40     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a373_1 ( .OUT(na373_1), .IN1(1'b1), .IN2(~na26_2), .IN3(1'b0), .IN4(1'b0), .IN5(na76_1), .IN6(na190_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x26y43     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a374_1 ( .OUT(na374_1), .IN1(1'b1), .IN2(na26_2), .IN3(1'b0), .IN4(1'b0), .IN5(na90_1), .IN6(na77_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x15y42     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a375_1 ( .OUT(na375_1), .IN1(1'b1), .IN2(~na73_1), .IN3(1'b0), .IN4(1'b0), .IN5(na103_1), .IN6(na79_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y62     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a376_4 ( .OUT(na376_2), .IN1(1'b1), .IN2(na77_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a376_6 ( .RAM_O2(na376_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na376_2), .COMP_OUT(1'b0) );
// C_MX2b////      x11y39     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a377_1 ( .OUT(na377_1), .IN1(1'b1), .IN2(na26_2), .IN3(1'b0), .IN4(1'b0), .IN5(na192_1), .IN6(na483_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x20y33     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a378_1 ( .OUT(na378_1), .IN1(1'b1), .IN2(na26_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na131_2), .IN8(na197_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x17y40     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a379_1 ( .OUT(na379_1), .IN1(1'b1), .IN2(na26_2), .IN3(1'b0), .IN4(1'b0), .IN5(na192_2), .IN6(na482_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y62     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a380_1 ( .OUT(na380_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na96_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a380_6 ( .RAM_O1(na380_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na380_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x23y35     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a381_1 ( .OUT(na381_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na467_2), .IN5(na92_1), .IN6(1'b0), .IN7(na199_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x18y37     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a382_1 ( .OUT(na382_1), .IN1(1'b1), .IN2(~na26_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na199_1), .IN8(na93_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x18y32     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a383_1 ( .OUT(na383_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na467_2), .IN5(1'b0), .IN6(na94_1), .IN7(1'b0), .IN8(na201_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x19y47     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a384_1 ( .OUT(na384_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na468_2), .IN5(na96_1), .IN6(1'b0), .IN7(na29_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y61     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a385_4 ( .OUT(na385_2), .IN1(na96_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a385_6 ( .RAM_O2(na385_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na385_2), .COMP_OUT(1'b0) );
// C_MX2b////      x24y37     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a386_1 ( .OUT(na386_1), .IN1(1'b1), .IN2(na26_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na9_2), .IN8(na201_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y61     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a387_1 ( .OUT(na387_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na28_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a387_6 ( .RAM_O1(na387_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na387_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x22y34     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a388_1 ( .OUT(na388_1), .IN1(1'b1), .IN2(~na26_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na195_1), .IN8(na102_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x17y33     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a389_1 ( .OUT(na389_1), .IN1(1'b1), .IN2(~na26_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na195_2), .IN8(na102_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y60     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a390_4 ( .OUT(na390_2), .IN1(1'b1), .IN2(na28_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a390_6 ( .RAM_O2(na390_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na390_2), .COMP_OUT(1'b0) );
// C_MX2b////      x20y43     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a391_1 ( .OUT(na391_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na468_2), .IN5(na76_1), .IN6(1'b0), .IN7(na486_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a392_1 ( .OUT(na392_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a392_6 ( .RAM_O1(na392_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na392_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x14y41     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a393_1 ( .OUT(na393_1), .IN1(na37_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na125_1), .IN8(na60_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y59     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a394_4 ( .OUT(na394_2), .IN1(1'b1), .IN2(1'b1), .IN3(na23_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a394_6 ( .RAM_O2(na394_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na394_2), .COMP_OUT(1'b0) );
// C_MX2b////      x24y42     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a395_1 ( .OUT(na395_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na468_2), .IN5(1'b0), .IN6(na28_2), .IN7(1'b0), .IN8(na27_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x22y33     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a396_1 ( .OUT(na396_1), .IN1(1'b1), .IN2(na26_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na131_1), .IN8(na197_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y59     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a397_1 ( .OUT(na397_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na24_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a397_6 ( .RAM_O1(na397_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na397_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y58     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a398_4 ( .OUT(na398_2), .IN1(1'b1), .IN2(1'b1), .IN3(na23_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a398_6 ( .RAM_O2(na398_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na398_2), .COMP_OUT(1'b0) );
// C_AND////      x28y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a399_1 ( .OUT(na399_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a399_6 ( .RAM_O1(na399_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na399_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a400_4 ( .OUT(na400_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a400_6 ( .RAM_O2(na400_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na400_2), .COMP_OUT(1'b0) );
// C_///AND/      x18y43     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a401_4 ( .OUT(na401_2), .IN1(na138_1), .IN2(na115_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x20y41     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a402_1 ( .OUT(na402_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na475_2), .IN6(1'b1), .IN7(~na39_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x1y95     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a403_4 ( .OUT(na403_2), .IN1(na67_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a403_6 ( .RAM_O2(na403_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na403_2), .COMP_OUT(1'b0) );
// C_///AND/      x19y1     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a404_4 ( .OUT(na404_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na141_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a404_6 ( .RAM_O2(na404_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na404_2), .COMP_OUT(1'b0) );
// C_AND////      x28y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a405_1 ( .OUT(na405_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a405_6 ( .RAM_O1(na405_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na405_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a406_4 ( .OUT(na406_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a406_6 ( .RAM_O2(na406_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na406_2), .COMP_OUT(1'b0) );
// C_AND////      x37y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a407_1 ( .OUT(na407_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a407_6 ( .RAM_O1(na407_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na407_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a408_4 ( .OUT(na408_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a408_6 ( .RAM_O2(na408_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na408_2), .COMP_OUT(1'b0) );
// C_AND////      x37y63     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a409_1 ( .OUT(na409_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na124_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a409_6 ( .RAM_O1(na409_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na409_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y62     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a410_4 ( .OUT(na410_2), .IN1(1'b1), .IN2(1'b1), .IN3(na123_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a410_6 ( .RAM_O2(na410_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na410_2), .COMP_OUT(1'b0) );
// C_AND////      x37y62     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a411_1 ( .OUT(na411_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na122_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a411_6 ( .RAM_O1(na411_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na411_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y61     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a412_4 ( .OUT(na412_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na121_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a412_6 ( .RAM_O2(na412_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na412_2), .COMP_OUT(1'b0) );
// C_AND////      x37y61     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a413_1 ( .OUT(na413_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na120_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a413_6 ( .RAM_O1(na413_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na413_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y60     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a414_4 ( .OUT(na414_2), .IN1(1'b1), .IN2(1'b1), .IN3(na119_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a414_6 ( .RAM_O2(na414_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na414_2), .COMP_OUT(1'b0) );
// C_AND////      x37y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a415_1 ( .OUT(na415_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a415_6 ( .RAM_O1(na415_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na415_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y59     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a416_4 ( .OUT(na416_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na118_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a416_6 ( .RAM_O2(na416_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na416_2), .COMP_OUT(1'b0) );
// C_AND////      x37y59     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a417_1 ( .OUT(na417_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na117_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a417_6 ( .RAM_O1(na417_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na417_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y58     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a418_4 ( .OUT(na418_2), .IN1(1'b1), .IN2(1'b1), .IN3(na116_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a418_6 ( .RAM_O2(na418_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na418_2), .COMP_OUT(1'b0) );
// C_AND////      x37y58     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a419_1 ( .OUT(na419_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a419_6 ( .RAM_O1(na419_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na419_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y57     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a420_4 ( .OUT(na420_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a420_6 ( .RAM_O2(na420_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na420_2), .COMP_OUT(1'b0) );
// C_AND////      x37y57     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a421_1 ( .OUT(na421_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a421_6 ( .RAM_O1(na421_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na421_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a422_4 ( .OUT(na422_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a422_6 ( .RAM_O2(na422_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na422_2), .COMP_OUT(1'b0) );
// C_AND////      x30y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a423_1 ( .OUT(na423_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a423_6 ( .RAM_O1(na423_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na423_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a424_4 ( .OUT(na424_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a424_6 ( .RAM_O2(na424_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na424_2), .COMP_OUT(1'b0) );
// C_AND////      x30y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a425_1 ( .OUT(na425_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a425_6 ( .RAM_O1(na425_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na425_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a426_4 ( .OUT(na426_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a426_6 ( .RAM_O2(na426_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na426_2), .COMP_OUT(1'b0) );
// C_AND////      x32y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a427_1 ( .OUT(na427_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a427_6 ( .RAM_O1(na427_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na427_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a428_4 ( .OUT(na428_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a428_6 ( .RAM_O2(na428_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na428_2), .COMP_OUT(1'b0) );
// C_AND////      x32y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a429_1 ( .OUT(na429_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a429_6 ( .RAM_O1(na429_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na429_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y62     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a430_4 ( .OUT(na430_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a430_6 ( .RAM_O2(na430_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na430_2), .COMP_OUT(1'b0) );
// C_AND////      x32y62     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a431_1 ( .OUT(na431_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a431_6 ( .RAM_O1(na431_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na431_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y61     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a432_4 ( .OUT(na432_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a432_6 ( .RAM_O2(na432_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na432_2), .COMP_OUT(1'b0) );
// C_AND////      x32y61     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a433_1 ( .OUT(na433_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a433_6 ( .RAM_O1(na433_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na433_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y60     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a434_4 ( .OUT(na434_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a434_6 ( .RAM_O2(na434_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na434_2), .COMP_OUT(1'b0) );
// C_AND////      x32y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a435_1 ( .OUT(na435_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a435_6 ( .RAM_O1(na435_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na435_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y59     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a436_4 ( .OUT(na436_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a436_6 ( .RAM_O2(na436_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na436_2), .COMP_OUT(1'b0) );
// C_AND////      x32y59     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a437_1 ( .OUT(na437_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na333_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a437_6 ( .RAM_O1(na437_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na437_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y58     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a438_4 ( .OUT(na438_2), .IN1(1'b1), .IN2(na205_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a438_6 ( .RAM_O2(na438_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na438_2), .COMP_OUT(1'b0) );
// C_AND////      x32y58     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a439_1 ( .OUT(na439_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na346_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a439_6 ( .RAM_O1(na439_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na439_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y57     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a440_4 ( .OUT(na440_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na345_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a440_6 ( .RAM_O2(na440_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na440_2), .COMP_OUT(1'b0) );
// C_AND////      x32y57     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a441_1 ( .OUT(na441_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na113_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a441_6 ( .RAM_O1(na441_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na441_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a442_4 ( .OUT(na442_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a442_6 ( .RAM_O2(na442_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na442_2), .COMP_OUT(1'b0) );
// C_AND////      x29y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a443_1 ( .OUT(na443_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a443_6 ( .RAM_O1(na443_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na443_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a444_4 ( .OUT(na444_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a444_6 ( .RAM_O2(na444_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na444_2), .COMP_OUT(1'b0) );
// C_AND////      x29y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a445_1 ( .OUT(na445_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a445_6 ( .RAM_O1(na445_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na445_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y64     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a446_4 ( .OUT(na446_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a446_6 ( .RAM_O2(na446_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na446_2), .COMP_OUT(1'b0) );
// C_AND////      x31y64     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a447_1 ( .OUT(na447_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a447_6 ( .RAM_O1(na447_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na447_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y63     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a448_4 ( .OUT(na448_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a448_6 ( .RAM_O2(na448_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na448_2), .COMP_OUT(1'b0) );
// C_AND////      x31y63     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a449_1 ( .OUT(na449_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a449_6 ( .RAM_O1(na449_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na449_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y62     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a450_4 ( .OUT(na450_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a450_6 ( .RAM_O2(na450_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na450_2), .COMP_OUT(1'b0) );
// C_AND////      x31y62     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a451_1 ( .OUT(na451_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a451_6 ( .RAM_O1(na451_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na451_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y61     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a452_4 ( .OUT(na452_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a452_6 ( .RAM_O2(na452_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na452_2), .COMP_OUT(1'b0) );
// C_AND////      x31y61     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a453_1 ( .OUT(na453_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a453_6 ( .RAM_O1(na453_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na453_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y60     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a454_4 ( .OUT(na454_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a454_6 ( .RAM_O2(na454_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na454_2), .COMP_OUT(1'b0) );
// C_AND////      x31y60     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a455_1 ( .OUT(na455_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a455_6 ( .RAM_O1(na455_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na455_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y59     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a456_4 ( .OUT(na456_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CINX(1'b0),
                     .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a456_6 ( .RAM_O2(na456_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na456_2), .COMP_OUT(1'b0) );
// C_/RAM_I1///      x34y59     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a457_2 ( .OUT(na457_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na341_96), .CP_O(1'b0) );
// C_////RAM_I2      x34y58     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a458_5 ( .OUT(na458_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na341_97), .CP_O(1'b0) );
// C_/RAM_I1///      x34y58     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a459_2 ( .OUT(na459_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na341_98), .CP_O(1'b0) );
// C_////RAM_I2      x34y57     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a460_5 ( .OUT(na460_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na341_99), .CP_O(1'b0) );
// C_/RAM_I1///      x34y57     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a461_2 ( .OUT(na461_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na341_100), .CP_O(1'b0) );
// C_////Bridge      x20y27     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a462_5 ( .OUT(na462_2), .IN1(na2_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y34     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a463_5 ( .OUT(na463_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na14_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y33     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a464_5 ( .OUT(na464_2), .IN1(na14_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x18y37     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a465_5 ( .OUT(na465_2), .IN1(na14_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x15y45     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a466_5 ( .OUT(na466_2), .IN1(1'b0), .IN2(1'b0), .IN3(na23_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y32     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a467_5 ( .OUT(na467_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na26_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y42     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a468_5 ( .OUT(na468_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na26_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x15y34     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a469_5 ( .OUT(na469_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na27_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y40     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a470_5 ( .OUT(na470_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na27_2) );
// C_////Bridge      x16y38     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a471_5 ( .OUT(na471_2), .IN1(1'b0), .IN2(1'b0), .IN3(na29_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y37     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a472_5 ( .OUT(na472_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na31_2) );
// C_////Bridge      x26y44     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a473_5 ( .OUT(na473_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na33_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y49     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a474_5 ( .OUT(na474_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na36_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y41     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a475_5 ( .OUT(na475_2), .IN1(1'b0), .IN2(1'b0), .IN3(na39_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x11y40     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a476_5 ( .OUT(na476_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na55_2) );
// C_////Bridge      x25y43     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a477_5 ( .OUT(na477_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na58_2), .IN8(1'b0) );
// C_////Bridge      x15y35     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a478_5 ( .OUT(na478_2), .IN1(1'b0), .IN2(1'b0), .IN3(na62_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y37     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a479_5 ( .OUT(na479_2), .IN1(1'b0), .IN2(1'b0), .IN3(na62_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x16y47     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a480_5 ( .OUT(na480_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na75_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y36     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a481_5 ( .OUT(na481_2), .IN1(na76_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y40     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a482_5 ( .OUT(na482_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na90_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x13y40     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a483_5 ( .OUT(na483_2), .IN1(na90_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y39     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a484_5 ( .OUT(na484_2), .IN1(1'b0), .IN2(na91_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y40     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a485_5 ( .OUT(na485_2), .IN1(1'b0), .IN2(na91_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y45     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a486_5 ( .OUT(na486_2), .IN1(na96_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y29     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a487_5 ( .OUT(na487_2), .IN1(1'b0), .IN2(1'b0), .IN3(na100_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y42     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a488_5 ( .OUT(na488_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na108_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x16y40     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a489_5 ( .OUT(na489_2), .IN1(1'b0), .IN2(na115_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y35     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a490_5 ( .OUT(na490_2), .IN1(1'b0), .IN2(na115_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y48     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a491_5 ( .OUT(na491_2), .IN1(1'b0), .IN2(1'b0), .IN3(na116_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x15y44     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a492_5 ( .OUT(na492_2), .IN1(na126_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y33     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a493_5 ( .OUT(na493_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na139_2) );
// C_////Bridge      x20y46     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a494_5 ( .OUT(na494_2), .IN1(1'b0), .IN2(1'b0), .IN3(na168_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y44     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a495_5 ( .OUT(na495_2), .IN1(1'b0), .IN2(1'b0), .IN3(na168_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x18y44     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a496_5 ( .OUT(na496_2), .IN1(1'b0), .IN2(1'b0), .IN3(na172_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y48     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a497_5 ( .OUT(na497_2), .IN1(1'b0), .IN2(1'b0), .IN3(na172_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y47     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a498_5 ( .OUT(na498_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na179_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y43     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a499_5 ( .OUT(na499_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na179_2) );
// C_////Bridge      x24y47     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a500_5 ( .OUT(na500_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na183_1) );
// C_////Bridge      x26y43     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a501_5 ( .OUT(na501_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na183_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
endmodule
