//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 July 2024)
//  Compile Time: 2024-07-19 12:30:06
//  Program Run:  2024-07-22 19:31:17
//  Program Call: /home/tibrahimovic/0.git-repo/cc-toolchain-linux/cc-toolchain-linux/bin/p_r/p_r -i net/top_synth.v -o top -ccf /home/tibrahimovic/projects/2.Simple--1/3.build/../1.hw/constraints/constraints.ccf -cCP --verbose 
//  File Type:    Verilog

// Gatecount:    510
module top (arst_n , clk , uart_rx ,
       led , o_psram_csn , o_psram_sclk , sent , tick_1us , uart_tx ,
       io_psram_data0 , io_psram_data1 , io_psram_data2 , io_psram_data3 , io_psram_data4 , io_psram_data5 , 
       io_psram_data6 , io_psram_data7 
) ;

input  arst_n;
input  clk;
input  uart_rx;

output led;
output o_psram_csn;
output o_psram_sclk;
output sent;
output tick_1us;
output uart_tx;

inout  io_psram_data0;
inout  io_psram_data1;
inout  io_psram_data2;
inout  io_psram_data3;
inout  io_psram_data4;
inout  io_psram_data5;
inout  io_psram_data6;
inout  io_psram_data7;


wire clk;
wire led;
wire sent;
wire na1_1;
wire na2_1;
wire na3_1;
wire na4_1;
wire na5_2;
wire na6_1;
wire na8_1;
wire arst_n;
wire na10_2;
wire na11_1;
wire na11_1_i;
wire na12_1;
wire na14_1;
wire na16_1;
wire na17_2;
wire na18_1;
wire na20_1;
wire na21_2;
wire na23_1;
wire na25_1;
wire na26_1;
wire na26_1_i;
wire na26_2;
wire na26_2_i;
wire na27_1;
wire na28_1;
wire na28_1_i;
wire na29_1;
wire na30_1;
wire na30_1_i;
wire na30_2;
wire na30_2_i;
wire na31_1;
wire na31_2;
wire na33_1;
wire na33_1_i;
wire na33_2;
wire na33_2_i;
wire na34_1;
wire na34_1_i;
wire na36_2;
wire na36_2_i;
wire na38_2;
wire na38_2_i;
wire na39_1;
wire na39_1_i;
wire na39_2;
wire na39_2_i;
wire na41_2;
wire na41_2_i;
wire na42_1;
wire na42_2;
wire na45_1;
wire na46_1;
wire na49_1;
wire na49_2;
wire na53_1;
wire na53_1_i;
wire na53_2;
wire na53_2_i;
wire na55_1;
wire na56_1;
wire na56_1_i;
wire na58_2;
wire na60_2;
wire na60_2_i;
wire na61_1;
wire na62_1;
wire na62_2;
wire na63_1;
wire na64_1;
wire na64_1_i;
wire na64_2;
wire na64_2_i;
wire na65_1;
wire na65_1_i;
wire na66_2;
wire na66_2_i;
wire na67_1;
wire na67_1_i;
wire na68_1;
wire na68_1_i;
wire na69_2;
wire na69_2_i;
wire na70_2;
wire na70_2_i;
wire na71_2;
wire na71_2_i;
wire na72_1;
wire na72_1_i;
wire na73_1;
wire na73_1_i;
wire na74_1;
wire na74_1_i;
wire na75_2;
wire na75_2_i;
wire na76_2;
wire na76_2_i;
wire na77_2;
wire na77_2_i;
wire na78_1;
wire na78_1_i;
wire na79_1;
wire na79_1_i;
wire na80_1;
wire na80_1_i;
wire na81_2;
wire na81_2_i;
wire na82_1;
wire na82_1_i;
wire na86_1;
wire na86_2;
wire na88_1;
wire na89_1;
wire na89_1_i;
wire na89_2;
wire na89_2_i;
wire na90_2;
wire na90_2_i;
wire na92_2;
wire na92_2_i;
wire na93_1;
wire na93_1_i;
wire na96_1;
wire na96_1_i;
wire na97_1;
wire na97_2;
wire na98_1;
wire na98_1_i;
wire na99_1;
wire na99_1_i;
wire na100_1;
wire na100_1_i;
wire na101_1;
wire na101_1_i;
wire na102_1;
wire na102_1_i;
wire na103_1;
wire na103_1_i;
wire na104_1;
wire na104_1_i;
wire na105_1;
wire na105_1_i;
wire na106_2;
wire na107_2;
wire na107_2_i;
wire na108_1;
wire na108_1_i;
wire na110_1;
wire na110_2;
wire na111_1;
wire na111_2;
wire na112_1;
wire na114_1;
wire na114_2;
wire na115_1;
wire na117_1;
wire na117_2;
wire na118_2;
wire na119_1;
wire na120_1;
wire na121_1;
wire na123_1;
wire na123_2;
wire na125_1;
wire na127_1;
wire na128_1;
wire na130_1;
wire na130_2;
wire na133_2;
wire na135_1;
wire na136_1;
wire na136_2;
wire na137_2;
wire na138_1;
wire na139_1;
wire na140_1;
wire na141_1;
wire na141_1_i;
wire na142_1;
wire na144_1;
wire na144_2;
wire na146_2;
wire na147_1;
wire na147_2;
wire na148_1;
wire na148_2;
wire na150_1;
wire na150_2;
wire na153_2;
wire na154_1;
wire na155_1;
wire na156_2;
wire na157_1;
wire na161_1;
wire na161_1_i;
wire na164_1;
wire na164_1_i;
wire na167_1;
wire na167_1_i;
wire na168_1;
wire na169_1;
wire na169_1_i;
wire na171_1;
wire na171_2;
wire na173_1;
wire na173_2;
wire na175_1;
wire na178_1;
wire na179_1;
wire na180_1;
wire na182_1;
wire na182_1_i;
wire na186_1;
wire na186_2;
wire na187_2;
wire na188_1;
wire na190_1;
wire na192_1;
wire na192_1_i;
wire na199_1;
wire na199_1_i;
wire na202_2;
wire na203_1;
wire na205_2;
wire na206_2;
wire na208_1;
wire na208_1_i;
wire na210_1;
wire na210_1_i;
wire na212_1;
wire na212_1_i;
wire na214_1;
wire na214_1_i;
wire na216_1;
wire na216_2;
wire na218_1;
wire na219_2;
wire na220_1;
wire na221_2;
wire na221_2_i;
wire na224_2;
wire na225_1;
wire na225_1_i;
wire na226_1;
wire na226_2;
wire na227_1;
wire na228_2;
wire na230_2;
wire na231_2;
wire na232_1;
wire na234_1;
wire na234_1_i;
wire na235_2;
wire na235_2_i;
wire na236_2;
wire na237_1;
wire na237_1_i;
wire na238_1;
wire na238_1_i;
wire na240_1;
wire na242_2;
wire na245_2;
wire na249_1;
wire na255_1;
wire na257_1;
wire na258_1;
wire na258_1_i;
wire na259_1;
wire na262_2;
wire na265_1;
wire na266_1;
wire na266_2;
wire na267_1;
wire na268_1;
wire na269_2;
wire na270_1;
wire na271_1;
wire na272_2;
wire na276_1;
wire na277_1;
wire na278_1;
wire na279_1;
wire na280_1;
wire na280_2;
wire na281_1;
wire na282_1;
wire na283_1;
wire na284_1;
wire na285_1;
wire na286_1;
wire na287_1;
wire na288_1;
wire na288_1_i;
wire na289_1;
wire na293_1;
wire na295_1;
wire na295_1_i;
wire na296_2;
wire na297_1;
wire na299_1;
wire na299_2;
wire na301_1;
wire na301_4;
wire na303_1;
wire na303_1_i;
wire na303_2;
wire na303_4;
wire na305_1;
wire na305_1_i;
wire na305_2;
wire na305_4;
wire na307_1;
wire na307_1_i;
wire na307_2;
wire na307_4;
wire na309_1;
wire na309_1_i;
wire na309_2;
wire na309_4;
wire na311_1;
wire na311_1_i;
wire na311_2;
wire na311_4;
wire na312_1;
wire na312_1_i;
wire na312_2;
wire na312_4;
wire na314_1;
wire na314_1_i;
wire na314_2;
wire na314_4;
wire na316_1;
wire na316_1_i;
wire na316_2;
wire na316_4;
wire na318_1;
wire na318_1_i;
wire na318_2;
wire na318_4;
wire na320_1;
wire na320_1_i;
wire na322_1;
wire na322_1_i;
wire na322_2;
wire na322_4;
wire na324_1;
wire na324_1_i;
wire na324_2;
wire na324_4;
wire na326_1;
wire na326_1_i;
wire na326_2;
wire na326_4;
wire na328_1;
wire na328_1_i;
wire na328_2;
wire na328_4;
wire na329_1;
wire na329_4;
wire na330_1;
wire na330_2;
wire na332_1;
wire na332_4;
wire na333_1;
wire na333_2;
wire na333_4;
wire na335_1;
wire na335_2;
wire na335_4;
wire na337_1;
wire na338_1;
wire na338_4;
wire na339_1;
wire na339_2;
wire na339_4;
wire na341_1;
wire na342_1;
wire na342_4;
wire na344_1;
wire na344_1_i;
wire na344_2;
wire na344_4;
wire na346_1;
wire na346_1_i;
wire na346_2;
wire na348_1;
wire na348_1_i;
wire na348_2;
wire na348_4;
wire na350_1;
wire na350_1_i;
wire na350_2;
wire na350_4;
wire na352_1;
wire na352_1_i;
wire na352_2;
wire na352_4;
wire na354_1;
wire na354_1_i;
wire na354_2;
wire na354_4;
wire na356_1;
wire na356_1_i;
wire na356_2;
wire na356_4;
wire na357_1;
wire na357_4;
wire na358_1;
wire na358_2;
wire na358_4;
wire na360_1;
wire na361_1;
wire na361_4;
wire na362_1;
wire na362_2;
wire na362_4;
wire na364_1;
wire na366_1;
wire na366_1_i;
wire na367_1;
wire na368_2;
wire na368_2_i;
wire na370_1;
wire na370_1_i;
wire na370_2;
wire na370_2_i;
wire na374_1;
wire na374_1_i;
wire na374_2;
wire na374_2_i;
wire na375_1;
wire na375_1_i;
wire na375_2;
wire na375_2_i;
wire na376_1;
wire na376_1_i;
wire na376_2;
wire na376_2_i;
wire na378_2;
wire na378_2_i;
wire na382_2;
wire na382_2_i;
wire na385_1;
wire na385_1_i;
wire na385_2;
wire na385_2_i;
wire na387_1;
wire na387_1_i;
wire na389_2;
wire na389_2_i;
wire na391_1;
wire na391_1_i;
wire na393_1;
wire na393_1_i;
wire na395_1;
wire na395_1_i;
wire na397_2;
wire na397_2_i;
wire na399_1;
wire na399_1_i;
wire na401_2;
wire na401_2_i;
wire na403_1;
wire na403_1_i;
wire na405_1;
wire na405_1_i;
wire na407_1;
wire na407_1_i;
wire na409_2;
wire na409_2_i;
wire na430_1;
wire na430_1_i;
wire na438_1;
wire na438_1_i;
wire na438_2;
wire na438_2_i;
wire na442_1;
wire na442_1_i;
wire na442_2;
wire na442_2_i;
wire na443_1;
wire na443_1_i;
wire na443_2;
wire na443_2_i;
wire na444_1;
wire na444_1_i;
wire na444_2;
wire na444_2_i;
wire na446_2;
wire na446_2_i;
wire na447_2;
wire na447_2_i;
wire na448_2;
wire na448_2_i;
wire na449_1;
wire na449_1_i;
wire na450_2;
wire na450_2_i;
wire na451_1;
wire na451_1_i;
wire na452_2;
wire na452_2_i;
wire na453_2;
wire na453_2_i;
wire na454_2;
wire na454_2_i;
wire na455_1;
wire na455_1_i;
wire na456_2;
wire na456_2_i;
wire na457_1;
wire na457_1_i;
wire na458_1;
wire na458_1_i;
wire na459_1;
wire na459_1_i;
wire na460_2;
wire na460_2_i;
wire na461_1;
wire na461_1_i;
wire na462_2;
wire na462_2_i;
wire na463_1;
wire na463_1_i;
wire na463_2;
wire na463_2_i;
wire na464_1;
wire na464_1_i;
wire na465_1;
wire na465_1_i;
wire na465_2;
wire na465_2_i;
wire na466_1;
wire na466_1_i;
wire na468_1;
wire na468_1_i;
wire na470_2;
wire na470_2_i;
wire na471_1;
wire na471_1_i;
wire na472_2;
wire na472_2_i;
wire na473_2;
wire na473_2_i;
wire na474_2;
wire na474_2_i;
wire na475_1;
wire na475_1_i;
wire na476_2;
wire na476_2_i;
wire na477_1;
wire na477_1_i;
wire na484_2;
wire na484_2_i;
wire na485_2;
wire na485_2_i;
wire na486_2;
wire na486_2_i;
wire na487_1;
wire na487_1_i;
wire na488_2;
wire na488_2_i;
wire na489_1;
wire na489_1_i;
wire na490_1;
wire na490_1_i;
wire na491_1;
wire na491_1_i;
wire na492_2;
wire na492_2_i;
wire na493_1;
wire na493_1_i;
wire na494_2;
wire na494_2_i;
wire na497_1;
wire na497_1_i;
wire na500_1;
wire na500_1_i;
wire na501_1;
wire na501_1_i;
wire na501_2;
wire na501_2_i;
wire na502_1;
wire na502_1_i;
wire na502_2;
wire na502_2_i;
wire na503_1;
wire na503_1_i;
wire na504_2;
wire na504_2_i;
wire na532_1;
wire na532_1_i;
wire na532_2;
wire na532_2_i;
wire na533_1;
wire na533_1_i;
wire na533_2;
wire na533_2_i;
wire na534_1;
wire na534_1_i;
wire na534_2;
wire na534_2_i;
wire na538_1;
wire na538_1_i;
wire na538_2;
wire na538_2_i;
wire na539_1;
wire na539_1_i;
wire na540_2;
wire na540_2_i;
wire na542_1;
wire na542_1_i;
wire na542_2;
wire na542_2_i;
wire na543_2;
wire na543_2_i;
wire na546_1;
wire na546_1_i;
wire na546_2;
wire na546_2_i;
wire na547_2;
wire na547_2_i;
wire na548_1;
wire na548_1_i;
wire na550_1;
wire na550_1_i;
wire na550_2;
wire na550_2_i;
wire na556_2;
wire na556_2_i;
wire na567_1;
wire na567_1_i;
wire na567_2;
wire na567_2_i;
wire na569_1;
wire na569_1_i;
wire na573_2;
wire na573_2_i;
wire na575_2;
wire na575_2_i;
wire na577_1;
wire na577_1_i;
wire na577_2;
wire na577_2_i;
wire na579_2;
wire na579_2_i;
wire na581_1;
wire na581_1_i;
wire na582_2;
wire na582_2_i;
wire na583_1;
wire na583_1_i;
wire na584_1;
wire na584_1_i;
wire na585_1;
wire na585_1_i;
wire na586_2;
wire na586_2_i;
wire na587_1;
wire na587_1_i;
wire na588_2;
wire na588_2_i;
wire na590_1;
wire na590_1_i;
wire na591_1;
wire na591_1_i;
wire na592_1;
wire na592_1_i;
wire na593_2;
wire na593_2_i;
wire na594_1;
wire na594_1_i;
wire na595_2;
wire na595_2_i;
wire na596_2;
wire na596_2_i;
wire na597_2;
wire na597_2_i;
wire na598_1;
wire na598_1_i;
wire na600_1;
wire na601_1;
wire na602_1;
wire na603_1;
wire na604_1;
wire na605_1;
wire na606_1;
wire na607_1;
wire na608_1;
wire na609_1;
wire na610_1;
wire na611_1;
wire na617_1;
wire na619_1;
wire na620_2;
wire na620_2_i;
wire na621_1;
wire na621_4;
wire na622_1;
wire na624_1;
wire na625_1;
wire na629_1;
wire na630_2;
wire na631_1;
wire na633_1;
wire na634_1;
wire na639_1;
wire na644_1;
wire na650_2;
wire na651_1;
wire na651_2;
wire na652_1;
wire na655_1;
wire na656_2;
wire na660_1;
wire na667_1;
wire na671_1;
wire na679_1;
wire na680_2;
wire na681_2;
wire na683_1;
wire na683_2;
wire na685_1;
wire na686_1;
wire na694_2;
wire na695_1;
wire na696_1;
wire na697_1;
wire na698_1;
wire na698_2;
wire na702_2;
wire na703_1;
wire na703_2;
wire na704_1;
wire na705_1;
wire na705_2;
wire na706_1;
wire na706_2;
wire na710_1;
wire na710_2;
wire na711_2;
wire na713_2;
wire na714_1;
wire na715_1;
wire na716_1;
wire na716_2;
wire na718_2;
wire na719_1;
wire na720_2;
wire na721_1;
wire na723_1;
wire na724_2;
wire na726_1;
wire na727_1;
wire na729_2;
wire na730_2;
wire na736_2;
wire na737_1;
wire na737_2;
wire na746_2;
wire na752_1;
wire na752_2;
wire na753_1;
wire na755_1;
wire na757_1;
wire na758_1;
wire na759_2;
wire na762_1;
wire na765_1;
wire na766_2;
wire na767_2;
wire na768_2;
wire na769_2;
wire na770_2;
wire na771_2;
wire na772_2;
wire na773_2;
wire na774_2;
wire na775_2;
wire na776_2;
wire na777_2;
wire na778_2;
wire na779_2;
wire na780_2;
wire na781_2;
wire na782_2;
wire na783_2;
wire na784_2;
wire na785_2;
wire na786_2;
wire na787_2;
wire na788_2;
wire na789_2;
wire na790_2;
wire na791_2;
wire na792_2;
wire na793_2;
wire na794_2;
wire na795_2;
wire na796_2;
wire na797_2;
wire na798_2;
wire na799_2;
wire na800_2;
wire na801_2;
wire na802_2;
wire na803_2;
wire na804_2;
wire na805_2;
wire na806_2;
wire na807_2;
wire na808_2;
wire na809_2;
wire na810_2;
wire na811_2;
wire na812_2;
wire na813_2;
wire na814_2;
wire na815_2;
wire na816_2;
wire na817_2;
wire na818_2;
wire na819_2;
wire na820_2;
wire na821_2;
wire na822_2;
wire na823_2;
wire na824_2;
wire na825_2;
wire na826_2;
wire na827_2;
wire na828_2;
wire na829_2;
wire na830_2;
wire na831_2;
wire na832_2;
wire na833_2;
wire na834_2;
wire na835_2;
wire na836_2;
wire na837_2;
wire na838_2;
wire na839_2;
wire na840_2;
wire na841_2;
wire na842_2;
wire na843_2;
wire na844_2;
wire na845_2;
wire na846_2;
wire na847_2;
wire na848_2;
wire na849_2;
wire na850_2;
wire na851_2;
wire na852_2;
wire uart_rx;
wire uart_tx;
wire na766_10;
wire na767_10;
wire na768_10;
wire na769_10;
wire na770_10;
wire na771_10;
wire na772_10;
wire na773_10;
wire na774_10;
wire na775_10;
wire na776_10;
wire na777_10;
wire na778_10;
wire na779_10;
wire na780_10;
wire na781_10;
wire na782_10;
wire na783_10;
wire na784_10;
wire na785_10;
wire na786_10;
wire na787_10;
wire tick_1us;
wire o_psram_csn;
wire o_psram_sclk;
wire io_psram_data0;
wire io_psram_data1;
wire io_psram_data2;
wire io_psram_data3;
wire io_psram_data4;
wire io_psram_data5;
wire io_psram_data6;
wire io_psram_data7;

// C_OR////      x101y30     80'h00_0018_00_0000_0CEE_0B00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1_1 ( .OUT(na1_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na619_1), .IN6(~na602_1), .IN7(1'b0), .IN8(1'b0),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x104y25     80'h00_0018_00_0000_0888_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2_1 ( .OUT(na2_1), .IN1(~na438_1), .IN2(~na442_1), .IN3(~na443_1), .IN4(~na444_1), .IN5(~na438_2), .IN6(~na442_2), .IN7(~na443_2),
                   .IN8(~na444_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a3 ( .PCLK0(na3_1), .PCLK1(_d0), .PCLK2(_d1), .PCLK3(_d2), .CLK0(na603_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0), .SER_CLK(1'b0),
                 .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_AND////      x107y23     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4_1 ( .OUT(na4_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na438_1), .IN6(~na848_2), .IN7(~na443_2), .IN8(~na444_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x100y26     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5_4 ( .OUT(na5_2), .IN1(1'b1), .IN2(~na1_1), .IN3(1'b1), .IN4(~na6_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x98y26     80'h00_0018_00_0000_0888_FEC5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a6_1 ( .OUT(na6_1), .IN1(~na543_2), .IN2(1'b0), .IN3(1'b0), .IN4(na752_2), .IN5(na66_2), .IN6(na93_1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x92y27     80'h00_0018_00_0000_0888_F151
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1), .IN1(~na542_2), .IN2(~na546_1), .IN3(~na547_2), .IN4(1'b1), .IN5(~na542_1), .IN6(~na546_2), .IN7(1'b1),
                   .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x93y21     80'h00_0060_00_0000_0C08_FF13
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a10_4 ( .OUT(na10_2), .IN1(1'b1), .IN2(~na548_1), .IN3(~na225_1), .IN4(~na550_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x100y8     80'h00_EE00_00_0000_0CEE_EC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a11_1 ( .OUT(na11_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na237_1), .IN7(na16_1), .IN8(na12_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a11_2 ( .OUT(na11_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na11_1_i) );
// C_AND////      x102y12     80'h00_0018_00_0000_0C88_4AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na622_1), .IN6(1'b1), .IN7(~na497_1), .IN8(na14_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y14     80'h00_0018_00_0000_0888_1F1C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a14_1 ( .OUT(na14_1), .IN1(1'b1), .IN2(na31_2), .IN3(~na26_1), .IN4(~na11_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na26_2), .IN8(~na28_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x96y7     80'h00_0018_00_0040_0C8C_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a16_1 ( .OUT(na16_1), .IN1(1'b0), .IN2(1'b0), .IN3(na789_2), .IN4(~na11_1), .IN5(1'b1), .IN6(na17_2), .IN7(1'b1), .IN8(~na790_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y8     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a17_4 ( .OUT(na17_2), .IN1(~na624_1), .IN2(na31_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x94y7     80'h00_0018_00_0000_0888_5153
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a18_1 ( .OUT(na18_1), .IN1(1'b1), .IN2(~na501_1), .IN3(~na502_2), .IN4(1'b1), .IN5(~na504_2), .IN6(~na501_2), .IN7(~na502_1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y10     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a20_1 ( .OUT(na20_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na849_2), .IN6(~na500_1), .IN7(~na221_2), .IN8(~na503_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x95y11     80'h00_0060_00_0000_0C08_FF45
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a21_4 ( .OUT(na21_2), .IN1(~na849_2), .IN2(1'b1), .IN3(~na18_1), .IN4(na14_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y13     80'h00_0018_00_0000_0C88_42FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a23_1 ( .OUT(na23_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na622_1), .IN6(~na237_1), .IN7(~na497_1), .IN8(na14_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x102y8     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a25_1 ( .OUT(na25_1), .IN1(1'b1), .IN2(na17_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na26_2), .IN8(~na362_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D//OR/D      x100y9     80'h00_EE00_80_0000_0CEE_CEAA
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a26_1 ( .OUT(na26_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na27_1), .IN6(na237_1), .IN7(1'b0), .IN8(na12_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a26_2 ( .OUT(na26_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na26_1_i) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a26_4 ( .OUT(na26_2_i), .IN1(na625_1), .IN2(1'b0), .IN3(na23_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a26_5 ( .OUT(na26_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na26_2_i) );
// C_MX4a////      x97y9     80'h00_0018_00_0040_0C0C_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1), .IN1(1'b0), .IN2(1'b0), .IN3(na26_1), .IN4(na362_2), .IN5(1'b1), .IN6(na17_2), .IN7(1'b1), .IN8(~na790_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x100y12     80'h00_EE00_00_0000_0788_F3E5
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a28_1 ( .OUT(na28_1_i), .IN1(~na21_2), .IN2(1'b0), .IN3(na29_1), .IN4(na12_1), .IN5(1'b0), .IN6(~na237_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a28_2 ( .OUT(na28_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na28_1_i) );
// C_MX2b////      x96y11     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a29_1 ( .OUT(na29_1), .IN1(1'b1), .IN2(~na17_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na364_1), .IN8(~na28_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x90y10     80'h00_EE00_80_0000_0C88_33A3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a30_1 ( .OUT(na30_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na31_1), .IN7(1'b1), .IN8(~na30_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a30_2 ( .OUT(na30_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na30_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a30_4 ( .OUT(na30_2_i), .IN1(1'b1), .IN2(~na31_1), .IN3(na335_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a30_5 ( .OUT(na30_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na30_2_i) );
// C_AND////D      x89y16     80'h00_FA18_00_0000_0888_4F41
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a31_1 ( .OUT(na31_1), .IN1(~na36_2), .IN2(~na34_1), .IN3(~na33_1), .IN4(na30_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na33_2),
                    .IN8(na30_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a31_5 ( .OUT(na31_2), .CLK(na367_1), .EN(na602_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na31_1) );
// C_AND/D//AND/D      x90y15     80'h00_EE00_80_0000_0C88_C3C3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_1 ( .OUT(na33_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na31_1), .IN7(1'b1), .IN8(na333_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_2 ( .OUT(na33_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na33_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a33_4 ( .OUT(na33_2_i), .IN1(1'b1), .IN2(~na31_1), .IN3(1'b1), .IN4(na337_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a33_5 ( .OUT(na33_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na33_2_i) );
// C_AND/D///      x89y10     80'h00_EE00_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a34_1 ( .OUT(na34_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na31_1), .IN7(1'b1), .IN8(na333_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a34_2 ( .OUT(na34_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na34_1_i) );
// C_///AND/D      x91y11     80'h00_EE00_80_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a36_4 ( .OUT(na36_2_i), .IN1(1'b1), .IN2(~na31_1), .IN3(na335_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a36_5 ( .OUT(na36_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na36_2_i) );
// C_///AND/D      x101y26     80'h00_EA00_80_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a38_4 ( .OUT(na38_2_i), .IN1(1'b1), .IN2(na238_1), .IN3(~na795_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a38_5 ( .OUT(na38_2), .CLK(na367_1), .EN(na257_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na38_2_i) );
// C_AND/D//AND/D      x110y24     80'h00_EA00_80_0000_0C88_F8F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_1 ( .OUT(na39_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na299_1), .IN6(na238_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_2 ( .OUT(na39_1), .CLK(na367_1), .EN(na257_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na39_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a39_4 ( .OUT(na39_2_i), .IN1(na299_2), .IN2(na238_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a39_5 ( .OUT(na39_2), .CLK(na367_1), .EN(na257_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na39_2_i) );
// C_///OR/D      x93y14     80'h00_EE00_80_0000_0C0E_FFAE
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a41_4 ( .OUT(na41_2_i), .IN1(na629_1), .IN2(na49_1), .IN3(na235_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a41_5 ( .OUT(na41_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na41_2_i) );
// C_AND///AND/      x93y11     80'h00_0078_00_0000_0C88_4CAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a42_1 ( .OUT(na42_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na41_2), .IN7(~na630_2), .IN8(na793_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a42_4 ( .OUT(na42_2), .IN1(na10_2), .IN2(1'b1), .IN3(na633_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y21     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na8_1), .IN8(~na550_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y20     80'h00_0018_00_0000_0888_515C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a46_1 ( .OUT(na46_1), .IN1(1'b1), .IN2(na31_2), .IN3(~na53_1), .IN4(1'b1), .IN5(~na56_1), .IN6(~na41_2), .IN7(~na53_2),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x95y14     80'h00_0078_00_0000_0C88_F458
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a49_1 ( .OUT(na49_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na10_2), .IN6(na46_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a49_4 ( .OUT(na49_2), .IN1(na358_1), .IN2(na31_2), .IN3(~na630_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x96y15     80'h00_EE00_80_0000_0C88_F135
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a53_1 ( .OUT(na53_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na42_2), .IN6(~na639_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a53_2 ( .OUT(na53_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na53_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a53_4 ( .OUT(na53_2_i), .IN1(~na42_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na634_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a53_5 ( .OUT(na53_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na53_2_i) );
// C_AND////      x92y9     80'h00_0018_00_0000_0C88_58FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na358_2), .IN6(na31_2), .IN7(~na630_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x97y17     80'h00_EE00_00_0000_0788_FB53
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a56_1 ( .OUT(na56_1_i), .IN1(1'b0), .IN2(~na644_1), .IN3(~na235_2), .IN4(1'b0), .IN5(na45_1), .IN6(~na46_1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a56_2 ( .OUT(na56_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na56_1_i) );
// C_///AND/      x92y11     80'h00_0060_00_0000_0C08_FF43
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a58_4 ( .OUT(na58_2), .IN1(1'b1), .IN2(~na360_1), .IN3(~na630_2), .IN4(na792_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x101y29     80'h00_FA00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a60_4 ( .OUT(na60_2_i), .IN1(1'b1), .IN2(na341_1), .IN3(1'b1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a60_5 ( .OUT(na60_2), .CLK(na367_1), .EN(na268_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na60_2_i) );
// C_AND////      x102y30     80'h00_0018_00_0000_0888_1AA3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a61_1 ( .OUT(na61_1), .IN1(1'b1), .IN2(~na295_1), .IN3(na62_1), .IN4(1'b1), .IN5(na141_1), .IN6(1'b1), .IN7(~na161_1), .IN8(~na108_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x100y21     80'h00_0078_00_0000_0C88_C511
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a62_1 ( .OUT(na62_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na167_1), .IN6(1'b1), .IN7(1'b1), .IN8(na164_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a62_4 ( .OUT(na62_2), .IN1(~na141_1), .IN2(~na295_1), .IN3(~na161_1), .IN4(~na108_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y21     80'h00_0018_00_0000_0C88_12FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a63_1 ( .OUT(na63_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na141_1), .IN6(~na295_1), .IN7(~na161_1), .IN8(~na108_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x104y31     80'h00_FA00_80_0000_0C88_CA4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a64_1 ( .OUT(na64_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na339_2), .IN6(1'b1), .IN7(1'b1), .IN8(na61_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a64_2 ( .OUT(na64_1), .CLK(na367_1), .EN(na268_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na64_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a64_4 ( .OUT(na64_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na64_2), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a64_5 ( .OUT(na64_2), .CLK(na367_1), .EN(na268_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na64_2_i) );
// C_AND/D///      x105y32     80'h00_FA00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a65_1 ( .OUT(na65_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na339_1), .IN6(1'b1), .IN7(1'b1), .IN8(na61_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a65_2 ( .OUT(na65_1), .CLK(na367_1), .EN(na268_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na65_1_i) );
// C_///ORAND/D      x99y29     80'h00_F600_80_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a66_4 ( .OUT(na66_2_i), .IN1(na650_2), .IN2(~na788_2), .IN3(na602_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a66_5 ( .OUT(na66_2), .CLK(na367_1), .EN(~na5_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na66_2_i) );
// C_AND/D///      x93y24     80'h00_FA00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_1 ( .OUT(na67_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na602_1), .IN8(na588_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_2 ( .OUT(na67_1), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na67_1_i) );
// C_AND/D///      x100y28     80'h00_FA00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a68_1 ( .OUT(na68_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na602_1), .IN8(na587_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a68_2 ( .OUT(na68_1), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na68_1_i) );
// C_///AND/D      x97y32     80'h00_FA00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a69_4 ( .OUT(na69_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na586_2), .IN4(na602_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a69_5 ( .OUT(na69_2), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na69_2_i) );
// C_///AND/D      x101y32     80'h00_FA00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a70_4 ( .OUT(na70_2_i), .IN1(1'b1), .IN2(na585_1), .IN3(na602_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a70_5 ( .OUT(na70_2), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na70_2_i) );
// C_///AND/D      x103y26     80'h00_FA00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a71_4 ( .OUT(na71_2_i), .IN1(na584_1), .IN2(1'b1), .IN3(na602_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a71_5 ( .OUT(na71_2), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na71_2_i) );
// C_AND/D///      x99y32     80'h00_FA00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a72_1 ( .OUT(na72_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na583_1), .IN8(na602_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a72_2 ( .OUT(na72_1), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na72_1_i) );
// C_AND/D///      x97y32     80'h00_FA00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a73_1 ( .OUT(na73_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na602_1), .IN8(na582_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a73_2 ( .OUT(na73_1), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na73_1_i) );
// C_AND/D///      x93y28     80'h00_FA00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a74_1 ( .OUT(na74_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na581_1), .IN7(1'b1), .IN8(na602_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a74_2 ( .OUT(na74_1), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na74_1_i) );
// C_///AND/D      x101y23     80'h00_FA00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a75_4 ( .OUT(na75_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na602_1), .IN4(na598_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a75_5 ( .OUT(na75_2), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na75_2_i) );
// C_///AND/D      x102y27     80'h00_FA00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a76_4 ( .OUT(na76_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na597_2), .IN4(na602_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a76_5 ( .OUT(na76_2), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na76_2_i) );
// C_///AND/D      x93y27     80'h00_FA00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a77_4 ( .OUT(na77_2_i), .IN1(na596_2), .IN2(1'b1), .IN3(na602_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a77_5 ( .OUT(na77_2), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na77_2_i) );
// C_AND/D///      x97y29     80'h00_FA00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na595_2), .IN6(1'b1), .IN7(1'b1), .IN8(na602_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_2 ( .OUT(na78_1), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_1_i) );
// C_AND/D///      x99y25     80'h00_FA00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a79_1 ( .OUT(na79_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na594_1), .IN8(na602_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a79_2 ( .OUT(na79_1), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na79_1_i) );
// C_AND/D///      x99y31     80'h00_FA00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na593_2), .IN8(na602_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_2 ( .OUT(na80_1), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na80_1_i) );
// C_///AND/D      x93y31     80'h00_FA00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a81_4 ( .OUT(na81_2_i), .IN1(na592_1), .IN2(1'b1), .IN3(na602_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a81_5 ( .OUT(na81_2), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na81_2_i) );
// C_OR/DST///      x91y32     80'h20_BA00_00_0000_0EEE_EDE7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a82_1 ( .OUT(na82_1_i), .IN1(~na88_1), .IN2(~na652_1), .IN3(na86_1), .IN4(na651_1), .IN5(~na656_2), .IN6(na655_1), .IN7(na86_2),
                    .IN8(na651_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'b1_0100_0000)) 
           _a82_2 ( .OUT(na82_1), .CLK(na367_1), .EN(na259_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na82_1_i) );
// C_AND///AND/      x92y29     80'h00_0078_00_0000_0C88_CAAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a86_1 ( .OUT(na86_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na542_2), .IN6(1'b1), .IN7(1'b1), .IN8(na102_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a86_4 ( .OUT(na86_2), .IN1(na542_1), .IN2(1'b1), .IN3(na99_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x95y29     80'h00_0018_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a88_1 ( .OUT(na88_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na105_1), .IN6(~na546_1), .IN7(~na101_1), .IN8(~na550_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x96y20     80'h00_FA00_80_0000_0C88_8F4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na330_2), .IN8(na660_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_2 ( .OUT(na89_1), .CLK(na367_1), .EN(na216_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a89_4 ( .OUT(na89_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na805_2), .IN4(na660_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a89_5 ( .OUT(na89_2), .CLK(na367_1), .EN(na216_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_2_i) );
// C_///AND/D      x89y20     80'h00_FA00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a90_4 ( .OUT(na90_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na330_1), .IN4(na660_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a90_5 ( .OUT(na90_2), .CLK(na367_1), .EN(na216_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na90_2_i) );
// C_///AND/D      x93y23     80'h00_FA00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a92_4 ( .OUT(na92_2_i), .IN1(na591_1), .IN2(1'b1), .IN3(na602_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a92_5 ( .OUT(na92_2), .CLK(na367_1), .EN(na1_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na92_2_i) );
// C_AND/D///      x97y28     80'h00_F600_00_0000_0888_CAA1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_1 ( .OUT(na93_1_i), .IN1(~na543_2), .IN2(~na93_1), .IN3(na602_1), .IN4(1'b1), .IN5(na66_2), .IN6(1'b1), .IN7(1'b1),
                    .IN8(na752_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_2 ( .OUT(na93_1), .CLK(na367_1), .EN(~na5_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na93_1_i) );
// C_MX2b/D///      x89y31     80'h00_FA00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a96_1 ( .OUT(na96_1_i), .IN1(1'b1), .IN2(~na844_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na601_1), .IN8(na600_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a96_2 ( .OUT(na96_1), .CLK(na367_1), .EN(na281_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na96_1_i) );
// C_AND////D      x105y17     80'h00_EE18_00_0000_0888_8FF5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a97_1 ( .OUT(na97_1), .IN1(~na97_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na497_1), .IN8(na14_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a97_5 ( .OUT(na97_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na97_1) );
// C_MX2a/D///      x93y25     80'h00_EA00_00_0040_0C03_0200
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a98_1 ( .OUT(na98_1_i), .IN1(na92_2), .IN2(na74_1), .IN3(1'b0), .IN4(1'b0), .IN5(na66_2), .IN6(~na93_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a98_2 ( .OUT(na98_1), .CLK(na367_1), .EN(na224_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na98_1_i) );
// C_MX2b/D///      x96y29     80'h00_EA00_00_0040_0A30_0002
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a99_1 ( .OUT(na99_1_i), .IN1(na66_2), .IN2(~na93_1), .IN3(1'b0), .IN4(1'b0), .IN5(na81_2), .IN6(na73_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a99_2 ( .OUT(na99_1), .CLK(na367_1), .EN(na224_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                    .D_IN(na99_1_i) );
// C_MX2a/D///      x97y31     80'h00_EA00_00_0040_0C03_0200
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a100_1 ( .OUT(na100_1_i), .IN1(na80_1), .IN2(na72_1), .IN3(1'b0), .IN4(1'b0), .IN5(na66_2), .IN6(~na93_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a100_2 ( .OUT(na100_1), .CLK(na367_1), .EN(na224_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na100_1_i) );
// C_MX2a/D///      x98y27     80'h00_EA00_00_0040_0C03_0200
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a101_1 ( .OUT(na101_1_i), .IN1(na79_1), .IN2(na71_2), .IN3(1'b0), .IN4(1'b0), .IN5(na66_2), .IN6(~na93_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a101_2 ( .OUT(na101_1), .CLK(na367_1), .EN(na224_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na101_1_i) );
// C_MX2b/D///      x96y30     80'h00_EA00_00_0040_0A30_0002
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a102_1 ( .OUT(na102_1_i), .IN1(na66_2), .IN2(~na93_1), .IN3(1'b0), .IN4(1'b0), .IN5(na78_1), .IN6(na70_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a102_2 ( .OUT(na102_1), .CLK(na367_1), .EN(na224_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na102_1_i) );
// C_MX2a/D///      x94y29     80'h00_EA00_00_0040_0C03_0200
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_1 ( .OUT(na103_1_i), .IN1(na77_2), .IN2(na69_2), .IN3(1'b0), .IN4(1'b0), .IN5(na66_2), .IN6(~na93_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_2 ( .OUT(na103_1), .CLK(na367_1), .EN(na224_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na103_1_i) );
// C_MX2a/D///      x97y27     80'h00_EA00_00_0040_0C0C_F200
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a104_1 ( .OUT(na104_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na76_2), .IN4(na68_1), .IN5(na66_2), .IN6(~na93_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a104_2 ( .OUT(na104_1), .CLK(na367_1), .EN(na224_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na104_1_i) );
// C_MX2b/D///      x95y25     80'h00_EA00_00_0040_0A30_0002
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a105_1 ( .OUT(na105_1_i), .IN1(na66_2), .IN2(~na93_1), .IN3(1'b0), .IN4(1'b0), .IN5(na75_2), .IN6(na67_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a105_2 ( .OUT(na105_1), .CLK(na367_1), .EN(na224_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na105_1_i) );
// C_///AND/      x89y8     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a106_4 ( .OUT(na106_2), .IN1(na367_1), .IN2(~na620_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x104y23     80'h00_FA00_80_0000_0C08_FF42
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a107_4 ( .OUT(na107_2_i), .IN1(na797_2), .IN2(~na38_2), .IN3(~na288_1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a107_5 ( .OUT(na107_2), .CLK(na367_1), .EN(na249_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na107_2_i) );
// C_ORAND*/D///      x98y22     80'h00_EA00_00_0000_0788_E55C
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a108_1 ( .OUT(na108_1_i), .IN1(1'b0), .IN2(na115_1), .IN3(~na123_1), .IN4(1'b0), .IN5(~na818_2), .IN6(1'b0), .IN7(na667_1),
                     .IN8(na108_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a108_2 ( .OUT(na108_1), .CLK(na367_1), .EN(na271_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na108_1_i) );
// C_AND///AND/      x101y15     80'h00_0078_00_0000_0C88_CC85
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a110_1 ( .OUT(na110_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na112_1), .IN7(1'b1), .IN8(na111_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a110_4 ( .OUT(na110_2), .IN1(~na141_1), .IN2(1'b1), .IN3(na123_1), .IN4(na833_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x98y14     80'h00_0078_00_0000_0C88_35AC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a111_1 ( .OUT(na111_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na167_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na164_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a111_4 ( .OUT(na111_2), .IN1(1'b1), .IN2(na737_2), .IN3(na62_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y18     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a112_1 ( .OUT(na112_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na141_1), .IN6(~na295_1), .IN7(na161_1), .IN8(~na108_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x99y16     80'h00_0078_00_0000_0C88_1488
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a114_1 ( .OUT(na114_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na141_1), .IN6(na295_1), .IN7(~na161_1), .IN8(~na108_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a114_4 ( .OUT(na114_2), .IN1(na141_1), .IN2(na295_1), .IN3(na161_1), .IN4(na108_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x101y20     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a115_1 ( .OUT(na115_1), .IN1(~na167_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na121_1), .IN8(~na119_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x95y19     80'h00_0078_00_0000_0C88_2818
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a117_1 ( .OUT(na117_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na141_1), .IN6(na295_1), .IN7(na161_1), .IN8(~na108_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a117_4 ( .OUT(na117_2), .IN1(na141_1), .IN2(na295_1), .IN3(~na161_1), .IN4(~na108_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y16     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a118_4 ( .OUT(na118_2), .IN1(1'b1), .IN2(1'b1), .IN3(na120_1), .IN4(na119_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y18     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a119_1 ( .OUT(na119_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na295_1), .IN7(1'b1), .IN8(~na108_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x100y15     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a120_1 ( .OUT(na120_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na167_1), .IN6(~na824_2), .IN7(na161_1), .IN8(na164_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x104y15     80'h00_0018_00_0000_0C88_2AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a121_1 ( .OUT(na121_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na167_1), .IN6(1'b1), .IN7(na62_2), .IN8(~na164_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x102y21     80'h00_0078_00_0000_0C88_415A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a123_1 ( .OUT(na123_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na167_1), .IN6(~na295_1), .IN7(~na806_2), .IN8(na164_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a123_4 ( .OUT(na123_2), .IN1(na110_1), .IN2(1'b1), .IN3(~na107_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y21     80'h00_0018_00_0000_0C88_85FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a125_1 ( .OUT(na125_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na141_1), .IN6(1'b1), .IN7(na161_1), .IN8(na111_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y23     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a127_1 ( .OUT(na127_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na112_1), .IN7(na62_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x96y23     80'h00_0018_00_0000_0888_5C2A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1), .IN1(na141_1), .IN2(1'b1), .IN3(na62_1), .IN4(~na108_1), .IN5(1'b1), .IN6(na295_1), .IN7(~na161_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x97y13     80'h00_0078_00_0000_0C88_828C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a130_1 ( .OUT(na130_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na141_1), .IN6(~na295_1), .IN7(na161_1), .IN8(na108_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a130_4 ( .OUT(na130_2), .IN1(1'b1), .IN2(na112_1), .IN3(na107_2), .IN4(na111_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x98y18     80'h00_0060_00_0000_0C08_FFCE
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a133_4 ( .OUT(na133_2), .IN1(na810_2), .IN2(na737_2), .IN3(1'b0), .IN4(na111_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x97y24     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a135_1 ( .OUT(na135_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na295_1), .IN7(1'b1), .IN8(na108_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x105y20     80'h00_0078_00_0000_0C88_423A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a136_1 ( .OUT(na136_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na141_1), .IN6(~na671_1), .IN7(~na161_1), .IN8(na111_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a136_4 ( .OUT(na136_2), .IN1(na125_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na108_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x97y23     80'h00_0060_00_0000_0C0E_FFAD
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a137_4 ( .OUT(na137_2), .IN1(~na141_1), .IN2(na671_1), .IN3(na161_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x97y25     80'h00_0018_00_0040_0C12_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(1'b1), .IN2(na671_1), .IN3(1'b0), .IN4(1'b0), .IN5(na125_1), .IN6(1'b1), .IN7(~na139_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x100y25     80'h00_0018_00_0000_0CEE_5700
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a139_1 ( .OUT(na139_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na140_1), .IN6(~na135_1), .IN7(~na62_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y17     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a140_1 ( .OUT(na140_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na141_1), .IN6(1'b1), .IN7(~na161_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x97y19     80'h00_EA00_00_0000_0EEE_5DEE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a141_1 ( .OUT(na141_1_i), .IN1(na142_1), .IN2(na144_1), .IN3(na123_2), .IN4(na148_1), .IN5(~na146_2), .IN6(na144_2), .IN7(~na156_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a141_2 ( .OUT(na141_1), .CLK(na367_1), .EN(na271_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na141_1_i) );
// C_AND////      x99y17     80'h00_0018_00_0000_0888_1244
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a142_1 ( .OUT(na142_1), .IN1(~na110_1), .IN2(na154_1), .IN3(~na123_1), .IN4(na147_1), .IN5(na146_2), .IN6(~na144_1), .IN7(~na850_2),
                     .IN8(~na147_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x95y18     80'h00_0078_00_0000_0C88_AEAE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a144_1 ( .OUT(na144_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na117_2), .IN6(na150_2), .IN7(na62_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a144_4 ( .OUT(na144_2), .IN1(na117_1), .IN2(na150_1), .IN3(na62_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x99y23     80'h00_0060_00_0000_0C0E_FF5D
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a146_4 ( .OUT(na146_2), .IN1(~na140_1), .IN2(na295_1), .IN3(~na62_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x98y16     80'h00_0078_00_0000_0C88_138F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a147_1 ( .OUT(na147_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na144_2), .IN7(~na829_2), .IN8(~na111_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a147_4 ( .OUT(na147_2), .IN1(1'b1), .IN2(1'b1), .IN3(na679_1), .IN4(na111_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x102y20     80'h00_0078_00_0000_0C88_AEAE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a148_1 ( .OUT(na148_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na130_1), .IN6(na112_1), .IN7(na62_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a148_4 ( .OUT(na148_2), .IN1(na814_2), .IN2(na135_1), .IN3(na120_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x99y20     80'h00_0078_00_0000_0C88_8444
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a150_1 ( .OUT(na150_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na141_1), .IN6(na295_1), .IN7(na161_1), .IN8(na108_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a150_4 ( .OUT(na150_2), .IN1(~na141_1), .IN2(na295_1), .IN3(~na161_1), .IN4(na108_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y22     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a153_4 ( .OUT(na153_2), .IN1(1'b1), .IN2(na295_1), .IN3(1'b1), .IN4(na108_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y24     80'h00_0018_00_0000_0C88_24FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a154_1 ( .OUT(na154_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na831_2), .IN6(na157_1), .IN7(na156_2), .IN8(~na133_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y26     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a155_1 ( .OUT(na155_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na62_2), .IN8(na111_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x102y17     80'h00_0060_00_0000_0C0E_FF3C
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a156_4 ( .OUT(na156_2), .IN1(1'b0), .IN2(na680_2), .IN3(1'b0), .IN4(~na111_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x101y18     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a157_1 ( .OUT(na157_1), .IN1(~na167_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na681_2), .IN6(~na114_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x100y19     80'h00_EA00_00_0000_0EEE_EECE
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a161_1 ( .OUT(na161_1_i), .IN1(na142_1), .IN2(na828_2), .IN3(1'b0), .IN4(na148_1), .IN5(na110_2), .IN6(na144_2), .IN7(na807_2),
                     .IN8(na148_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a161_2 ( .OUT(na161_1), .CLK(na367_1), .EN(na271_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na161_1_i) );
// C_OR/D///      x100y14     80'h00_EA00_00_0000_0EEE_EEE7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a164_1 ( .OUT(na164_1_i), .IN1(~na683_1), .IN2(~na827_2), .IN3(na123_1), .IN4(na111_2), .IN5(na683_2), .IN6(na144_1), .IN7(na826_2),
                     .IN8(na148_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a164_2 ( .OUT(na164_1), .CLK(na367_1), .EN(na271_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na164_1_i) );
// C_AND*/D///      x101y17     80'h00_EA00_00_0000_0388_1FFF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a167_1 ( .OUT(na167_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na168_1), .IN8(~na817_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a167_2 ( .OUT(na167_1), .CLK(na367_1), .EN(na271_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na167_1_i) );
// C_AND////      x108y15     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a168_1 ( .OUT(na168_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na114_2), .IN7(na62_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*/D///      x109y11     80'h00_EA00_00_0000_0788_C814
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a169_1 ( .OUT(na169_1_i), .IN1(~na695_1), .IN2(na175_1), .IN3(~na686_1), .IN4(~na171_1), .IN5(na694_2), .IN6(na685_1), .IN7(1'b1),
                     .IN8(na171_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a169_2 ( .OUT(na169_1), .CLK(na367_1), .EN(na297_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na169_1_i) );
// C_AND///AND/      x106y14     80'h00_0078_00_0000_0C88_F211
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a171_1 ( .OUT(na171_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na462_2), .IN6(~na186_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a171_4 ( .OUT(na171_2), .IN1(~na130_2), .IN2(~na180_1), .IN3(~na179_1), .IN4(~na178_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x100y17     80'h00_0078_00_0000_0C88_AE73
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a173_1 ( .OUT(na173_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na117_1), .IN6(na150_2), .IN7(na62_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a173_4 ( .OUT(na173_2), .IN1(1'b0), .IN2(~na808_2), .IN3(~na62_1), .IN4(~na809_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x103y12     80'h00_0018_00_0000_0888_F373
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a175_1 ( .OUT(na175_1), .IN1(1'b0), .IN2(~na136_1), .IN3(~na819_2), .IN4(~na111_1), .IN5(1'b0), .IN6(~na136_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x102y24     80'h00_0018_00_0000_0888_EFAA
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a178_1 ( .OUT(na178_1), .IN1(na458_1), .IN2(1'b0), .IN3(na62_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na62_2), .IN8(na830_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x104y21     80'h00_0018_00_0000_0888_FEAC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a179_1 ( .OUT(na179_1), .IN1(1'b0), .IN2(na450_2), .IN3(na62_1), .IN4(1'b0), .IN5(na130_1), .IN6(na114_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x103y16     80'h00_0018_00_0000_0888_FEAC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a180_1 ( .OUT(na180_1), .IN1(1'b0), .IN2(na454_2), .IN3(na62_1), .IN4(1'b0), .IN5(na851_2), .IN6(na112_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x107y7     80'h00_EA00_00_0000_0EEE_AAB7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_1 ( .OUT(na182_1_i), .IN1(~na696_1), .IN2(~na175_1), .IN3(na703_1), .IN4(~na702_2), .IN5(na110_1), .IN6(1'b0), .IN7(na703_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_2 ( .OUT(na182_1), .CLK(na367_1), .EN(na297_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na182_1_i) );
// C_ORAND///ORAND/      x103y18     80'h00_0078_00_0000_0C88_7777
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a186_1 ( .OUT(na186_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na816_2), .IN6(~na815_2), .IN7(~na812_2), .IN8(~na111_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a186_4 ( .OUT(na186_2), .IN1(~na816_2), .IN2(~na135_1), .IN3(~na813_2), .IN4(~na111_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x100y11     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a187_4 ( .OUT(na187_2), .IN1(na683_2), .IN2(na451_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y10     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a188_1 ( .OUT(na188_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na447_2), .IN6(1'b1), .IN7(na173_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x104y20     80'h00_0018_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a190_1 ( .OUT(na190_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na803_2), .IN6(na150_1), .IN7(na62_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x110y11     80'h00_EA00_00_0000_0EEE_C5D5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a192_1 ( .OUT(na192_1_i), .IN1(~na710_1), .IN2(1'b0), .IN3(~na704_1), .IN4(na713_2), .IN5(~na710_2), .IN6(1'b0), .IN7(1'b0),
                     .IN8(na711_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a192_2 ( .OUT(na192_1), .CLK(na367_1), .EN(na297_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na192_1_i) );
// C_OR/D///      x110y15     80'h00_EA00_00_0000_0EEE_BDEB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a199_1 ( .OUT(na199_1_i), .IN1(na719_1), .IN2(~na714_1), .IN3(na123_2), .IN4(na205_2), .IN5(~na718_2), .IN6(na136_2), .IN7(na822_2),
                     .IN8(~na206_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a199_2 ( .OUT(na199_1), .CLK(na367_1), .EN(na297_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na199_1_i) );
// C_///AND/      x100y23     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a202_4 ( .OUT(na202_2), .IN1(na683_2), .IN2(1'b1), .IN3(na453_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y28     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a203_1 ( .OUT(na203_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na449_1), .IN7(na173_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x110y22     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a205_4 ( .OUT(na205_2), .IN1(1'b1), .IN2(na461_1), .IN3(1'b1), .IN4(na190_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x102y18     80'h00_0060_00_0000_0C08_FF75
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a206_4 ( .OUT(na206_2), .IN1(~na110_2), .IN2(1'b0), .IN3(~na819_2), .IN4(~na111_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*/D///      x108y10     80'h00_EA00_00_0000_0788_841C
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a208_1 ( .OUT(na208_1_i), .IN1(1'b1), .IN2(na175_1), .IN3(~na686_1), .IN4(~na171_1), .IN5(~na721_1), .IN6(na685_1), .IN7(na720_2),
                     .IN8(na171_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a208_2 ( .OUT(na208_1), .CLK(na367_1), .EN(na297_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na208_1_i) );
// C_OR/D///      x103y7     80'h00_EA00_00_0000_0EEE_AAB7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a210_1 ( .OUT(na210_1_i), .IN1(~na696_1), .IN2(~na175_1), .IN3(na724_2), .IN4(~na723_1), .IN5(na110_1), .IN6(1'b0), .IN7(na703_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a210_2 ( .OUT(na210_1), .CLK(na367_1), .EN(na297_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na210_1_i) );
// C_OR/D///      x109y10     80'h00_EA00_00_0000_0EEE_D0D5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a212_1 ( .OUT(na212_1_i), .IN1(~na710_1), .IN2(1'b0), .IN3(~na704_1), .IN4(na727_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na726_1),
                     .IN8(na711_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a212_2 ( .OUT(na212_1), .CLK(na367_1), .EN(na297_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na212_1_i) );
// C_OR/D///      x108y16     80'h00_EA00_00_0000_0EEE_BDEB
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a214_1 ( .OUT(na214_1_i), .IN1(na730_2), .IN2(~na714_1), .IN3(na123_2), .IN4(na205_2), .IN5(~na729_2), .IN6(na136_2), .IN7(na822_2),
                     .IN8(~na206_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a214_2 ( .OUT(na214_1), .CLK(na367_1), .EN(na297_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na214_1_i) );
// C_ICOMP////D      x89y23     80'h00_F618_00_0000_0888_FF56
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a216_1 ( .OUT(na216_1), .IN1(~na382_2), .IN2(na82_1), .IN3(na835_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a216_5 ( .OUT(na216_2), .CLK(na367_1), .EN(~na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na216_1) );
// C_AND////      x96y25     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a218_1 ( .OUT(na218_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na220_1), .IN6(1'b1), .IN7(~na219_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x90y19     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a219_4 ( .OUT(na219_2), .IN1(na216_1), .IN2(na90_2), .IN3(na805_2), .IN4(na89_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x91y27     80'h00_0018_00_0000_0C88_84FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a220_1 ( .OUT(na220_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na216_1), .IN6(na847_2), .IN7(na318_1), .IN8(na320_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND*/D      x94y11     80'h00_EE00_80_0000_0C07_FFDB
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a221_4 ( .OUT(na221_2_i), .IN1(na617_1), .IN2(~na237_1), .IN3(~na221_2), .IN4(na14_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a221_5 ( .OUT(na221_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na221_2_i) );
// C_///AND/      x94y26     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a224_4 ( .OUT(na224_2), .IN1(1'b1), .IN2(1'b1), .IN3(na235_2), .IN4(na6_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x98y23     80'h00_EE00_00_0000_0388_3DFF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a225_1 ( .OUT(na225_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na836_2), .IN6(na46_1), .IN7(1'b0), .IN8(~na224_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a225_2 ( .OUT(na225_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na225_1_i) );
// C_OR////DST      x103y10     80'h20_BA18_00_0000_0EEE_50A0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a226_1 ( .OUT(na226_1), .IN1(1'b0), .IN2(1'b0), .IN3(na736_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na227_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'b1_0100_0000)) 
           _a226_5 ( .OUT(na226_2), .CLK(na367_1), .EN(na278_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na226_1) );
// C_MX4b////      x102y13     80'h00_0018_00_0040_0A3F_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a227_1 ( .OUT(na227_1), .IN1(1'b1), .IN2(~na737_2), .IN3(1'b1), .IN4(na164_1), .IN5(~na167_1), .IN6(~na737_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x100y13     80'h00_0060_00_0000_0C08_FF43
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a228_4 ( .OUT(na228_2), .IN1(1'b1), .IN2(~na237_1), .IN3(~na497_1), .IN4(na14_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x110y20     80'h00_0060_00_0000_0C08_FF42
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a230_4 ( .OUT(na230_2), .IN1(na231_2), .IN2(~na38_2), .IN3(~na796_2), .IN4(na39_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y25     80'h00_0060_00_0000_0C08_FFA8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a231_4 ( .OUT(na231_2), .IN1(na97_2), .IN2(na238_1), .IN3(na602_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x109y20     80'h00_0018_00_0000_0C88_48FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a232_1 ( .OUT(na232_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na231_2), .IN6(na38_2), .IN7(~na796_2), .IN8(na39_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x102y23     80'h00_EE00_00_0000_0388_75FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a234_1 ( .OUT(na234_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na842_2), .IN6(1'b0), .IN7(~na234_1), .IN8(~na280_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a234_2 ( .OUT(na234_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na234_1_i) );
// C_///ORAND*/DST      x94y19     80'h20_BE00_80_0000_0C07_FFD7
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a235_4 ( .OUT(na235_2_i), .IN1(~na543_2), .IN2(~na46_1), .IN3(~na235_2), .IN4(na6_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'b1_0100_0100)) 
           _a235_5 ( .OUT(na235_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na235_2_i) );
// C_///AND/      x106y24     80'h00_0060_00_0000_0C08_FF18
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a236_4 ( .OUT(na236_2), .IN1(na231_2), .IN2(na38_2), .IN3(~na798_2), .IN4(~na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/DST///      x93y16     80'h20_BE00_00_0000_0388_77FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a237_1 ( .OUT(na237_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na617_1), .IN6(~na237_1), .IN7(~na497_1),
                     .IN8(~na14_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'b1_0100_0000)) 
           _a237_2 ( .OUT(na237_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na237_1_i) );
// C_ORAND*/D///      x107y22     80'h00_EE00_00_0000_0388_BBFF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a238_1 ( .OUT(na238_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na617_1), .IN6(~na258_1), .IN7(na839_2), .IN8(~na838_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a238_2 ( .OUT(na238_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na238_1_i) );
// C_ORAND////      x109y23     80'h00_0018_00_0000_0888_CFE3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a240_1 ( .OUT(na240_1), .IN1(1'b0), .IN2(~na38_2), .IN3(na2_1), .IN4(na39_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b0), .IN8(na39_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x105y23     80'h00_0060_00_0000_0C08_FF22
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a242_4 ( .OUT(na242_2), .IN1(na231_2), .IN2(~na38_2), .IN3(na796_2), .IN4(~na39_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x108y21     80'h00_0060_00_0000_0C08_FF28
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a245_4 ( .OUT(na245_2), .IN1(na231_2), .IN2(na38_2), .IN3(na796_2), .IN4(~na39_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x106y17     80'h00_0018_00_0000_0888_FEAB
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a249_1 ( .OUT(na249_1), .IN1(na240_1), .IN2(~na238_1), .IN3(na602_1), .IN4(1'b0), .IN5(na842_2), .IN6(na238_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y25     80'h00_0018_00_0000_0C88_12FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a255_1 ( .OUT(na255_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na231_2), .IN6(~na38_2), .IN7(~na798_2), .IN8(~na39_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x106y20     80'h00_0018_00_0040_0A70_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a257_1 ( .OUT(na257_1), .IN1(1'b1), .IN2(~na238_1), .IN3(1'b1), .IN4(na617_1), .IN5(na97_2), .IN6(na258_1), .IN7(na746_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/DST///      x103y22     80'h20_BE00_00_0000_0388_D7FF
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a258_1 ( .OUT(na258_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na617_1), .IN6(~na258_1), .IN7(~na234_1),
                     .IN8(na280_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'b1_0100_0000)) 
           _a258_2 ( .OUT(na258_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na258_1_i) );
// C_ORAND////      x95y22     80'h00_0018_00_0000_0888_BEDE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a259_1 ( .OUT(na259_1), .IN1(na852_2), .IN2(na46_1), .IN3(~na225_1), .IN4(na793_2), .IN5(na45_1), .IN6(na46_1), .IN7(na235_2),
                     .IN8(~na752_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x97y11     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a262_4 ( .OUT(na262_2), .IN1(1'b1), .IN2(na150_2), .IN3(1'b1), .IN4(na111_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x105y10     80'h00_0018_00_0040_0A31_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a265_1 ( .OUT(na265_1), .IN1(na110_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na753_1), .IN6(na430_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////DST      x108y8     80'h20_BA18_00_0000_0888_AF73
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a266_1 ( .OUT(na266_1), .IN1(1'b0), .IN2(~na802_2), .IN3(~na811_2), .IN4(~na111_1), .IN5(1'b1), .IN6(1'b1), .IN7(na227_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'b1_0100_0000)) 
           _a266_5 ( .OUT(na266_2), .CLK(na367_1), .EN(na265_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na266_1) );
// C_MX2b////      x107y8     80'h00_0018_00_0040_0A31_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a267_1 ( .OUT(na267_1), .IN1(na110_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na840_2), .IN6(na430_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x101y31     80'h00_0018_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a268_1 ( .OUT(na268_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na269_2), .IN6(na755_1), .IN7(na602_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y25     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a269_4 ( .OUT(na269_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na270_1), .IN4(na61_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x102y29     80'h00_0018_00_0000_0C88_81FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a270_1 ( .OUT(na270_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na60_2), .IN6(~na65_1), .IN7(na64_1), .IN8(na804_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x101y22     80'h00_0018_00_0000_0888_FDB5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a271_1 ( .OUT(na271_1), .IN1(~na272_2), .IN2(1'b0), .IN3(na270_1), .IN4(~na61_1), .IN5(~na110_1), .IN6(na430_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x105y29     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a272_4 ( .OUT(na272_2), .IN1(1'b1), .IN2(1'b1), .IN3(na757_1), .IN4(na155_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x107y29     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a276_1 ( .OUT(na276_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na569_1), .IN6(na567_1), .IN7(na350_1), .IN8(na348_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y8     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a277_1 ( .OUT(na277_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na737_2), .IN7(1'b1), .IN8(na111_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x101y11     80'h00_0018_00_0040_0A31_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a278_1 ( .OUT(na278_1), .IN1(na110_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na759_2), .IN6(na430_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x99y15     80'h00_0018_00_0040_0A31_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a279_1 ( .OUT(na279_1), .IN1(na110_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na841_2), .IN6(na430_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////DST      x106y22     80'h20_BA18_00_0000_0888_FF73
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a280_1 ( .OUT(na280_1), .IN1(1'b0), .IN2(~na226_1), .IN3(~na811_2), .IN4(~na111_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'b1_0100_0000)) 
           _a280_5 ( .OUT(na280_2), .CLK(na367_1), .EN(na279_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na280_1) );
// C_AND////      x89y26     80'h00_0018_00_0000_0C88_A2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a281_1 ( .OUT(na281_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na216_2), .IN6(~na378_2), .IN7(na407_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y17     80'h00_0018_00_0000_0C88_12FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a282_1 ( .OUT(na282_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na216_1), .IN6(~na90_2), .IN7(~na805_2), .IN8(~na89_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y22     80'h00_0018_00_0000_0C88_42FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a283_1 ( .OUT(na283_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na216_1), .IN6(~na90_2), .IN7(~na805_2), .IN8(na89_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y24     80'h00_0018_00_0000_0C88_48FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_1 ( .OUT(na284_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na216_1), .IN6(na90_2), .IN7(~na805_2), .IN8(na89_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x89y20     80'h00_0018_00_0000_0C88_28FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a285_1 ( .OUT(na285_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na216_1), .IN6(na90_2), .IN7(na805_2), .IN8(~na89_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y19     80'h00_0018_00_0000_0C88_18FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a286_1 ( .OUT(na286_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na216_1), .IN6(na90_2), .IN7(~na805_2), .IN8(~na89_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x90y24     80'h00_0018_00_0000_0C88_82FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a287_1 ( .OUT(na287_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na216_1), .IN6(~na90_2), .IN7(na805_2), .IN8(na89_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x108y19     80'h00_EE00_00_0000_0888_C3EC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a288_1 ( .OUT(na288_1_i), .IN1(1'b0), .IN2(na238_1), .IN3(na2_1), .IN4(na39_1), .IN5(1'b0), .IN6(~na38_2), .IN7(1'b0), .IN8(na39_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a288_2 ( .OUT(na288_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na288_1_i) );
// C_AND////      x89y21     80'h00_0018_00_0000_0C88_22FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a289_1 ( .OUT(na289_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na216_1), .IN6(~na90_2), .IN7(na805_2), .IN8(~na89_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x99y13     80'h00_0018_00_0000_0CEE_EE00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a293_1 ( .OUT(na293_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na117_1), .IN6(na737_2), .IN7(na811_2), .IN8(na820_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x95y26     80'h00_EA00_00_0000_0EEE_CEA5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a295_1 ( .OUT(na295_1_i), .IN1(~na138_1), .IN2(1'b0), .IN3(na128_1), .IN4(1'b0), .IN5(na762_1), .IN6(na136_1), .IN7(1'b0),
                     .IN8(na148_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a295_2 ( .OUT(na295_1), .CLK(na367_1), .EN(na271_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na295_1_i) );
// C_///AND/      x97y15     80'h00_0060_00_0000_0C08_FF84
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a296_4 ( .OUT(na296_2), .IN1(~na262_2), .IN2(na186_2), .IN3(na173_2), .IN4(na206_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x107y12     80'h00_0018_00_0040_0A31_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a297_1 ( .OUT(na297_1), .IN1(na110_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na765_1), .IN6(na430_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x107y19     80'h00_0078_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a299_1 ( .OUT(na299_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na38_2), .IN7(1'b1), .IN8(na39_1),
                     .CINX(1'b0), .CINY1(na301_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a299_4 ( .OUT(na299_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na39_2), .IN5(1'b1), .IN6(na38_2), .IN7(1'b1), .IN8(na39_1),
                     .CINX(1'b0), .CINY1(na301_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x107y18     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a301_2 ( .OUT(na301_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a301_6 ( .COUTY1(na301_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na301_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x92y18     80'h00_EE60_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a303_1 ( .OUT(na303_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na303_1),
                     .CINX(1'b0), .CINY1(na328_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a303_2 ( .OUT(na303_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na303_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a303_4 ( .OUT(na303_2), .COUTY1(na303_4), .IN1(na395_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na303_1), .CINX(1'b0), .CINY1(na328_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x92y19     80'h00_EE60_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a305_1 ( .OUT(na305_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na305_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na303_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a305_2 ( .OUT(na305_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na305_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a305_4 ( .OUT(na305_2), .COUTY1(na305_4), .IN1(na397_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na305_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na303_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x92y20     80'h00_EE60_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a307_1 ( .OUT(na307_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na307_1),
                     .CINX(1'b0), .CINY1(na305_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a307_2 ( .OUT(na307_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na307_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a307_4 ( .OUT(na307_2), .COUTY1(na307_4), .IN1(na399_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na307_1), .CINX(1'b0), .CINY1(na305_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x92y21     80'h00_EE60_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a309_1 ( .OUT(na309_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na309_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na307_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a309_2 ( .OUT(na309_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na309_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a309_4 ( .OUT(na309_2), .COUTY1(na309_4), .IN1(na401_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na309_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na307_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x92y22     80'h00_EE60_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a311_1 ( .OUT(na311_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na311_1),
                     .CINX(1'b0), .CINY1(na309_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a311_2 ( .OUT(na311_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na311_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a311_4 ( .OUT(na311_2), .COUTY1(na311_4), .IN1(na403_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na311_1), .CINX(1'b0), .CINY1(na309_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x92y13     80'h00_EE60_00_0020_0C66_AA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a312_1 ( .OUT(na312_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na385_2), .IN6(1'b1), .IN7(na312_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na329_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a312_2 ( .OUT(na312_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na312_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a312_4 ( .OUT(na312_2), .COUTY1(na312_4), .IN1(na385_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na385_2), .IN6(1'b1), .IN7(na312_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na329_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x92y23     80'h00_EE60_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a314_1 ( .OUT(na314_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na314_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na311_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a314_2 ( .OUT(na314_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na314_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a314_4 ( .OUT(na314_2), .COUTY1(na314_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na405_1), .IN5(1'b0), .IN6(1'b0), .IN7(na314_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na311_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x92y24     80'h00_EE60_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a316_1 ( .OUT(na316_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na316_1),
                     .CINX(1'b0), .CINY1(na314_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a316_2 ( .OUT(na316_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na316_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a316_4 ( .OUT(na316_2), .COUTY1(na316_4), .IN1(1'b0), .IN2(1'b0), .IN3(na407_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na316_1), .CINX(1'b0), .CINY1(na314_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x92y25     80'h00_EE60_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a318_1 ( .OUT(na318_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na318_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na316_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a318_2 ( .OUT(na318_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na318_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a318_4 ( .OUT(na318_2), .COUTY1(na318_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na409_2), .IN5(1'b0), .IN6(1'b0), .IN7(na318_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na316_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF/D///      x92y26     80'h00_EE00_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a320_1 ( .OUT(na320_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na320_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na318_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a320_2 ( .OUT(na320_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na320_1_i) );
// C_ADDF2/D//ADDF2/      x92y14     80'h00_EE60_00_0020_0C66_C00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a322_1 ( .OUT(na322_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na322_1),
                     .CINX(1'b0), .CINY1(na312_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a322_2 ( .OUT(na322_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na322_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a322_4 ( .OUT(na322_2), .COUTY1(na322_4), .IN1(1'b1), .IN2(na387_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na322_1), .CINX(1'b0), .CINY1(na312_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x92y15     80'h00_EE60_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a324_1 ( .OUT(na324_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na324_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na322_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a324_2 ( .OUT(na324_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na324_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a324_4 ( .OUT(na324_2), .COUTY1(na324_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na389_2), .IN5(1'b0), .IN6(1'b0), .IN7(na324_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na322_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x92y16     80'h00_EE60_00_0020_0C66_C00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a326_1 ( .OUT(na326_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na326_1),
                     .CINX(1'b0), .CINY1(na324_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a326_2 ( .OUT(na326_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na326_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a326_4 ( .OUT(na326_2), .COUTY1(na326_4), .IN1(1'b1), .IN2(na391_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na326_1), .CINX(1'b0), .CINY1(na324_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x92y17     80'h00_EE60_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a328_1 ( .OUT(na328_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na328_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na326_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a328_2 ( .OUT(na328_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na328_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a328_4 ( .OUT(na328_2), .COUTY1(na328_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na393_1), .IN5(1'b0), .IN6(1'b0), .IN7(na328_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na326_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x92y12     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a329_2 ( .OUT(na329_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a329_6 ( .COUTY1(na329_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na329_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x90y17     80'h00_0078_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a330_1 ( .OUT(na330_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na90_2), .IN7(1'b1), .IN8(na89_2),
                     .CINX(1'b0), .CINY1(na332_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a330_4 ( .OUT(na330_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na89_1), .IN5(1'b1), .IN6(na90_2), .IN7(1'b1), .IN8(na89_2),
                     .CINX(1'b0), .CINY1(na332_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x90y16     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a332_2 ( .OUT(na332_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a332_6 ( .COUTY1(na332_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na332_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x90y12     80'h00_0078_00_0020_0C66_CA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a333_1 ( .OUT(na333_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na794_2), .IN6(1'b1), .IN7(1'b1), .IN8(na30_1),
                     .CINX(1'b0), .CINY1(na338_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a333_4 ( .OUT(na333_2), .COUTY1(na333_4), .IN1(1'b1), .IN2(na34_1), .IN3(1'b0), .IN4(1'b0), .IN5(na794_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na30_1), .CINX(1'b0), .CINY1(na338_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x90y13     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a335_1 ( .OUT(na335_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na30_2),
                     .CINX(1'b0), .CINY1(na333_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a335_4 ( .OUT(na335_2), .COUTY1(na335_4), .IN1(na36_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na30_2), .CINX(1'b0), .CINY1(na333_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x90y14     80'h00_0018_00_0010_0666_00A0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a337_1 ( .OUT(na337_1), .IN1(1'b0), .IN2(1'b0), .IN3(na33_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na335_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x90y11     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a338_2 ( .OUT(na338_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a338_6 ( .COUTY1(na338_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na338_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x103y29     80'h00_0078_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a339_1 ( .OUT(na339_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na65_1), .IN7(na64_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na342_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a339_4 ( .OUT(na339_2), .COUTY1(na339_4), .IN1(1'b0), .IN2(1'b0), .IN3(na64_1), .IN4(1'b1), .IN5(1'b1), .IN6(na65_1), .IN7(na64_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na342_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x103y30     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a341_1 ( .OUT(na341_1), .IN1(na60_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na339_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x103y28     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a342_2 ( .OUT(na342_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a342_6 ( .COUTY1(na342_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na342_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x108y29     80'h00_EA60_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a344_1 ( .OUT(na344_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na344_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na356_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a344_2 ( .OUT(na344_1), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na344_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a344_4 ( .OUT(na344_2), .COUTY1(na344_4), .IN1(1'b1), .IN2(na577_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na344_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na356_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x108y30     80'h00_EA60_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a346_1 ( .OUT(na346_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na346_1),
                     .CINX(1'b0), .CINY1(na344_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a346_2 ( .OUT(na346_1), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na346_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a346_4 ( .OUT(na346_2), .IN1(na579_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na346_1),
                     .CINX(1'b0), .CINY1(na344_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x108y24     80'h00_EA60_00_0020_0C66_CC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a348_1 ( .OUT(na348_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na567_2), .IN7(1'b1), .IN8(na348_1),
                     .CINX(1'b0), .CINY1(na357_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a348_2 ( .OUT(na348_1), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na348_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a348_4 ( .OUT(na348_2), .COUTY1(na348_4), .IN1(1'b1), .IN2(na567_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na567_2), .IN7(1'b1),
                     .IN8(na348_1), .CINX(1'b0), .CINY1(na357_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x108y25     80'h00_EA60_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a350_1 ( .OUT(na350_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na350_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na348_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a350_2 ( .OUT(na350_1), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na350_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a350_4 ( .OUT(na350_2), .COUTY1(na350_4), .IN1(na569_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na350_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na348_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x108y26     80'h00_EA60_00_0020_0C66_C00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a352_1 ( .OUT(na352_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na352_1),
                     .CINX(1'b0), .CINY1(na350_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a352_2 ( .OUT(na352_1), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na352_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a352_4 ( .OUT(na352_2), .COUTY1(na352_4), .IN1(1'b1), .IN2(na577_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na352_1), .CINX(1'b0), .CINY1(na350_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x108y27     80'h00_EA60_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a354_1 ( .OUT(na354_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na354_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na352_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a354_2 ( .OUT(na354_1), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na354_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a354_4 ( .OUT(na354_2), .COUTY1(na354_4), .IN1(na573_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na354_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na352_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x108y28     80'h00_EA60_00_0020_0C66_C0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a356_1 ( .OUT(na356_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na356_1),
                     .CINX(1'b0), .CINY1(na354_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a356_2 ( .OUT(na356_1), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na356_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a356_4 ( .OUT(na356_2), .COUTY1(na356_4), .IN1(1'b0), .IN2(1'b0), .IN3(na575_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na356_1), .CINX(1'b0), .CINY1(na354_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x108y23     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a357_2 ( .OUT(na357_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a357_6 ( .COUTY1(na357_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na357_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x91y15     80'h00_0078_00_0020_0C66_ACAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a358_1 ( .OUT(na358_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na41_2), .IN7(na53_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na361_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a358_4 ( .OUT(na358_2), .COUTY1(na358_4), .IN1(1'b1), .IN2(1'b1), .IN3(na53_1), .IN4(1'b1), .IN5(1'b1), .IN6(na41_2), .IN7(na53_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na361_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x91y16     80'h00_0018_00_0010_0666_00FA
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a360_1 ( .OUT(na360_1), .IN1(na56_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na358_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x91y14     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a361_2 ( .OUT(na361_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a361_6 ( .COUTY1(na361_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na361_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x98y10     80'h00_0078_00_0020_0C66_CAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a362_1 ( .OUT(na362_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na791_2), .IN6(1'b1), .IN7(1'b1), .IN8(na11_1),
                     .CINX(1'b0), .CINY1(na621_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a362_4 ( .OUT(na362_2), .COUTY1(na362_4), .IN1(1'b1), .IN2(1'b1), .IN3(na26_1), .IN4(1'b1), .IN5(na791_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na11_1), .CINX(1'b0), .CINY1(na621_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x98y11     80'h00_0018_00_0010_0666_00CF
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a364_1 ( .OUT(na364_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na28_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na362_4), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x90y28     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a366_1 ( .OUT(na366_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na82_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a366_2 ( .OUT(na366_1), .CLK(na367_1), .EN(na289_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na366_1_i) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0000_0010)) 
           _a367 ( .GLB0(na367_1), .GLB1(_d3), .GLB2(_d4), .GLB3(_d5), .CLK_FB0(_d6), .CLK_FB1(_d7), .CLK_FB2(_d8), .CLK_FB3(_d9),
                   .CLK0_0(1'b0), .CLK0_90(1'b0), .CLK0_180(1'b0), .CLK0_270(1'b0), .CLK0_BYP(na3_1), .CLK1_0(1'b0), .CLK1_90(1'b0),
                   .CLK1_180(1'b0), .CLK1_270(1'b0), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0), .CLK2_270(1'b0),
                   .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0), .USR_GLB0(1'b0),
                   .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0), .USR_FB3(1'b0) );
// C_///AND/D      x90y23     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a368_4 ( .OUT(na368_2_i), .IN1(1'b1), .IN2(na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a368_5 ( .OUT(na368_2), .CLK(na367_1), .EN(na282_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na368_2_i) );
// C_AND/D//AND/D      x101y12     80'h00_EA00_80_0000_0C88_FCCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a370_1 ( .OUT(na370_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na370_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a370_2 ( .OUT(na370_1), .CLK(na367_1), .EN(na228_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na370_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a370_4 ( .OUT(na370_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na375_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a370_5 ( .OUT(na370_2), .CLK(na367_1), .EN(na228_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na370_2_i) );
// C_AND/D//AND/D      x106y27     80'h00_EA00_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a374_1 ( .OUT(na374_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na375_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a374_2 ( .OUT(na374_1), .CLK(na367_1), .EN(na228_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na374_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a374_4 ( .OUT(na374_2_i), .IN1(na617_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a374_5 ( .OUT(na374_2), .CLK(na367_1), .EN(na228_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na374_2_i) );
// C_AND/D//AND/D      x108y20     80'h00_EA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a375_1 ( .OUT(na375_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na376_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a375_2 ( .OUT(na375_1), .CLK(na367_1), .EN(na228_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na375_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a375_4 ( .OUT(na375_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na376_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a375_5 ( .OUT(na375_2), .CLK(na367_1), .EN(na228_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na375_2_i) );
// C_AND/D//AND/D      x106y25     80'h00_EA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a376_1 ( .OUT(na376_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na374_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a376_2 ( .OUT(na376_1), .CLK(na367_1), .EN(na228_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na376_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a376_4 ( .OUT(na376_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na374_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a376_5 ( .OUT(na376_2), .CLK(na367_1), .EN(na228_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na376_2_i) );
// C_///AND/D      x89y24     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a378_4 ( .OUT(na378_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na407_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a378_5 ( .OUT(na378_2), .CLK(na367_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na378_2_i) );
// C_///AND/D      x89y21     80'h00_FE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a382_4 ( .OUT(na382_2_i), .IN1(1'b1), .IN2(na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a382_5 ( .OUT(na382_2), .CLK(na367_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na382_2_i) );
// C_AND/D//AND/D      x93y9     80'h00_EE00_80_0000_0C88_AFF5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a385_1 ( .OUT(na385_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na312_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a385_2 ( .OUT(na385_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na385_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a385_4 ( .OUT(na385_2_i), .IN1(~na385_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a385_5 ( .OUT(na385_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na385_2_i) );
// C_AND/D///      x93y10     80'h00_EE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a387_1 ( .OUT(na387_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na322_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a387_2 ( .OUT(na387_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na387_1_i) );
// C_///AND/D      x92y10     80'h00_EE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a389_4 ( .OUT(na389_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na324_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a389_5 ( .OUT(na389_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na389_2_i) );
// C_AND/D///      x93y12     80'h00_EE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a391_1 ( .OUT(na391_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na326_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a391_2 ( .OUT(na391_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na391_1_i) );
// C_AND/D///      x96y12     80'h00_EE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a393_1 ( .OUT(na393_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na328_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a393_2 ( .OUT(na393_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na393_1_i) );
// C_AND/D///      x93y15     80'h00_EE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a395_1 ( .OUT(na395_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na303_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a395_2 ( .OUT(na395_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na395_1_i) );
// C_///AND/D      x89y17     80'h00_EE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a397_4 ( .OUT(na397_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na305_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a397_5 ( .OUT(na397_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na397_2_i) );
// C_AND/D///      x93y17     80'h00_EE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a399_1 ( .OUT(na399_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na307_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a399_2 ( .OUT(na399_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na399_1_i) );
// C_///AND/D      x93y17     80'h00_EE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a401_4 ( .OUT(na401_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na309_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a401_5 ( .OUT(na401_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na401_2_i) );
// C_AND/D///      x93y21     80'h00_EE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a403_1 ( .OUT(na403_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na311_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a403_2 ( .OUT(na403_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na403_1_i) );
// C_AND/D///      x94y22     80'h00_EE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a405_1 ( .OUT(na405_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na314_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a405_2 ( .OUT(na405_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na405_1_i) );
// C_AND/D///      x90y25     80'h00_EE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a407_1 ( .OUT(na407_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na316_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a407_2 ( .OUT(na407_1), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na407_1_i) );
// C_///AND/D      x90y22     80'h00_EE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a409_4 ( .OUT(na409_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na318_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a409_5 ( .OUT(na409_2), .CLK(na367_1), .EN(1'b1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na409_2_i) );
// C_AND/D///      x105y14     80'h00_FA00_00_0000_0C88_5FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a430_1 ( .OUT(na430_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na288_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a430_2 ( .OUT(na430_1), .CLK(na367_1), .EN(na249_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na430_1_i) );
// C_AND/D//AND/D      x105y21     80'h00_FA00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a438_1 ( .OUT(na438_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na532_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a438_2 ( .OUT(na438_1), .CLK(na367_1), .EN(na255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na438_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a438_4 ( .OUT(na438_2_i), .IN1(na532_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a438_5 ( .OUT(na438_2), .CLK(na367_1), .EN(na255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na438_2_i) );
// C_AND/D//AND/D      x105y30     80'h00_FA00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a442_1 ( .OUT(na442_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na538_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a442_2 ( .OUT(na442_1), .CLK(na367_1), .EN(na255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na442_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a442_4 ( .OUT(na442_2_i), .IN1(na538_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a442_5 ( .OUT(na442_2), .CLK(na367_1), .EN(na255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na442_2_i) );
// C_AND/D//AND/D      x106y21     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a443_1 ( .OUT(na443_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na533_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a443_2 ( .OUT(na443_1), .CLK(na367_1), .EN(na255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na443_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a443_4 ( .OUT(na443_2_i), .IN1(1'b1), .IN2(na533_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a443_5 ( .OUT(na443_2), .CLK(na367_1), .EN(na255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na443_2_i) );
// C_AND/D//AND/D      x104y26     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a444_1 ( .OUT(na444_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na534_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a444_2 ( .OUT(na444_1), .CLK(na367_1), .EN(na255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na444_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a444_4 ( .OUT(na444_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na534_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a444_5 ( .OUT(na444_2), .CLK(na367_1), .EN(na255_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na444_2_i) );
// C_///AND/D      x103y9     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a446_4 ( .OUT(na446_2_i), .IN1(na532_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a446_5 ( .OUT(na446_2), .CLK(na367_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na446_2_i) );
// C_///AND/D      x101y9     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a447_4 ( .OUT(na447_2_i), .IN1(na532_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a447_5 ( .OUT(na447_2), .CLK(na367_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na447_2_i) );
// C_///AND/D      x103y15     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a448_4 ( .OUT(na448_2_i), .IN1(1'b1), .IN2(na533_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a448_5 ( .OUT(na448_2), .CLK(na367_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na448_2_i) );
// C_AND/D///      x105y28     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a449_1 ( .OUT(na449_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na534_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a449_2 ( .OUT(na449_1), .CLK(na367_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na449_1_i) );
// C_///AND/D      x101y30     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a450_4 ( .OUT(na450_2_i), .IN1(na538_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a450_5 ( .OUT(na450_2), .CLK(na367_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na450_2_i) );
// C_AND/D///      x103y14     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a451_1 ( .OUT(na451_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na533_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a451_2 ( .OUT(na451_1), .CLK(na367_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na451_1_i) );
// C_///AND/D      x102y28     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a452_4 ( .OUT(na452_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a452_5 ( .OUT(na452_2), .CLK(na367_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na452_2_i) );
// C_///AND/D      x102y33     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a453_4 ( .OUT(na453_2_i), .IN1(na538_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a453_5 ( .OUT(na453_2), .CLK(na367_1), .EN(na236_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na453_2_i) );
// C_///AND/D      x101y10     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a454_4 ( .OUT(na454_2_i), .IN1(na532_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a454_5 ( .OUT(na454_2), .CLK(na367_1), .EN(na242_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na454_2_i) );
// C_AND/D///      x102y10     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a455_1 ( .OUT(na455_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na532_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a455_2 ( .OUT(na455_1), .CLK(na367_1), .EN(na242_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na455_1_i) );
// C_///AND/D      x106y16     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a456_4 ( .OUT(na456_2_i), .IN1(1'b1), .IN2(na533_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a456_5 ( .OUT(na456_2), .CLK(na367_1), .EN(na242_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na456_2_i) );
// C_AND/D///      x104y28     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a457_1 ( .OUT(na457_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na534_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a457_2 ( .OUT(na457_1), .CLK(na367_1), .EN(na242_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na457_1_i) );
// C_AND/D///      x101y27     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a458_1 ( .OUT(na458_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na538_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a458_2 ( .OUT(na458_1), .CLK(na367_1), .EN(na242_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na458_1_i) );
// C_AND/D///      x108y13     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a459_1 ( .OUT(na459_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na533_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a459_2 ( .OUT(na459_1), .CLK(na367_1), .EN(na242_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na459_1_i) );
// C_///AND/D      x111y23     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a460_4 ( .OUT(na460_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a460_5 ( .OUT(na460_2), .CLK(na367_1), .EN(na242_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na460_2_i) );
// C_AND/D///      x105y26     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a461_1 ( .OUT(na461_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na538_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a461_2 ( .OUT(na461_1), .CLK(na367_1), .EN(na242_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na461_1_i) );
// C_///AND/D      x105y13     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a462_4 ( .OUT(na462_2_i), .IN1(na532_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a462_5 ( .OUT(na462_2), .CLK(na367_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na462_2_i) );
// C_AND/D//AND/D      x104y12     80'h00_FA00_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a463_1 ( .OUT(na463_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na532_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a463_2 ( .OUT(na463_1), .CLK(na367_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na463_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a463_4 ( .OUT(na463_2_i), .IN1(1'b1), .IN2(na533_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a463_5 ( .OUT(na463_2), .CLK(na367_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na463_2_i) );
// C_AND/D///      x107y17     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a464_1 ( .OUT(na464_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na533_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a464_2 ( .OUT(na464_1), .CLK(na367_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na464_1_i) );
// C_AND/D//AND/D      x105y31     80'h00_FA00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a465_1 ( .OUT(na465_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na534_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a465_2 ( .OUT(na465_1), .CLK(na367_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na465_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a465_4 ( .OUT(na465_2_i), .IN1(na538_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a465_5 ( .OUT(na465_2), .CLK(na367_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na465_2_i) );
// C_AND/D///      x109y21     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a466_1 ( .OUT(na466_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na538_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a466_2 ( .OUT(na466_1), .CLK(na367_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na466_1_i) );
// C_AND/D///      x110y20     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a468_1 ( .OUT(na468_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na534_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a468_2 ( .OUT(na468_1), .CLK(na367_1), .EN(na245_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na468_1_i) );
// C_///AND/D      x105y9     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a470_4 ( .OUT(na470_2_i), .IN1(na532_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a470_5 ( .OUT(na470_2), .CLK(na367_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na470_2_i) );
// C_AND/D///      x105y9     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a471_1 ( .OUT(na471_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na532_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a471_2 ( .OUT(na471_1), .CLK(na367_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na471_1_i) );
// C_///AND/D      x107y16     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a472_4 ( .OUT(na472_2_i), .IN1(1'b1), .IN2(na533_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a472_5 ( .OUT(na472_2), .CLK(na367_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na472_2_i) );
// C_///AND/D      x105y25     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a473_4 ( .OUT(na473_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na534_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a473_5 ( .OUT(na473_2), .CLK(na367_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na473_2_i) );
// C_///AND/D      x104y27     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a474_4 ( .OUT(na474_2_i), .IN1(na538_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a474_5 ( .OUT(na474_2), .CLK(na367_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na474_2_i) );
// C_AND/D///      x107y16     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a475_1 ( .OUT(na475_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na533_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a475_2 ( .OUT(na475_1), .CLK(na367_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na475_1_i) );
// C_///AND/D      x112y24     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a476_4 ( .OUT(na476_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na534_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a476_5 ( .OUT(na476_2), .CLK(na367_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na476_2_i) );
// C_AND/D///      x107y28     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a477_1 ( .OUT(na477_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na538_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a477_2 ( .OUT(na477_1), .CLK(na367_1), .EN(na230_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na477_1_i) );
// C_///AND/D      x106y10     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a484_4 ( .OUT(na484_2_i), .IN1(na532_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a484_5 ( .OUT(na484_2), .CLK(na367_1), .EN(na232_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na484_2_i) );
// C_///AND/D      x109y7     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a485_4 ( .OUT(na485_2_i), .IN1(na532_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a485_5 ( .OUT(na485_2), .CLK(na367_1), .EN(na232_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na485_2_i) );
// C_///AND/D      x107y13     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a486_4 ( .OUT(na486_2_i), .IN1(1'b1), .IN2(na533_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a486_5 ( .OUT(na486_2), .CLK(na367_1), .EN(na232_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na486_2_i) );
// C_AND/D///      x112y23     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a487_1 ( .OUT(na487_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na534_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a487_2 ( .OUT(na487_1), .CLK(na367_1), .EN(na232_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na487_1_i) );
// C_///AND/D      x106y28     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a488_4 ( .OUT(na488_2_i), .IN1(na538_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a488_5 ( .OUT(na488_2), .CLK(na367_1), .EN(na232_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na488_2_i) );
// C_AND/D///      x107y13     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a489_1 ( .OUT(na489_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na533_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a489_2 ( .OUT(na489_1), .CLK(na367_1), .EN(na232_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na489_1_i) );
// C_AND/D///      x109y22     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a490_1 ( .OUT(na490_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na534_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a490_2 ( .OUT(na490_1), .CLK(na367_1), .EN(na232_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na490_1_i) );
// C_AND/D///      x107y26     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a491_1 ( .OUT(na491_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na538_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a491_2 ( .OUT(na491_1), .CLK(na367_1), .EN(na232_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na491_1_i) );
// C_///AND/D      x91y28     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a492_4 ( .OUT(na492_2_i), .IN1(1'b1), .IN2(na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a492_5 ( .OUT(na492_2), .CLK(na367_1), .EN(na284_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na492_2_i) );
// C_AND/D///      x90y27     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a493_1 ( .OUT(na493_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na82_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a493_2 ( .OUT(na493_1), .CLK(na367_1), .EN(na287_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na493_1_i) );
// C_///AND/D      x91y31     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a494_4 ( .OUT(na494_2_i), .IN1(1'b1), .IN2(na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a494_5 ( .OUT(na494_2), .CLK(na367_1), .EN(na219_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na494_2_i) );
// C_AND/D///      x98y15     80'h00_EA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a497_1 ( .OUT(na497_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na504_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a497_2 ( .OUT(na497_1), .CLK(na367_1), .EN(na14_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na497_1_i) );
// C_AND/D///      x97y8     80'h00_EA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a500_1 ( .OUT(na500_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na502_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a500_2 ( .OUT(na500_1), .CLK(na367_1), .EN(na14_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na500_1_i) );
// C_AND/D//AND/D      x95y10     80'h00_EA00_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a501_1 ( .OUT(na501_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na221_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a501_2 ( .OUT(na501_1), .CLK(na367_1), .EN(na14_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na501_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a501_4 ( .OUT(na501_2_i), .IN1(1'b1), .IN2(na501_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a501_5 ( .OUT(na501_2), .CLK(na367_1), .EN(na14_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na501_2_i) );
// C_AND/D//AND/D      x92y7     80'h00_EA00_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a502_1 ( .OUT(na502_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na502_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a502_2 ( .OUT(na502_1), .CLK(na367_1), .EN(na14_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na502_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a502_4 ( .OUT(na502_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na503_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a502_5 ( .OUT(na502_2), .CLK(na367_1), .EN(na14_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na502_2_i) );
// C_AND/D///      x96y10     80'h00_EA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a503_1 ( .OUT(na503_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na501_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a503_2 ( .OUT(na503_1), .CLK(na367_1), .EN(na14_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na503_1_i) );
// C_///AND/D      x91y9     80'h00_EA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a504_4 ( .OUT(na504_2_i), .IN1(1'b1), .IN2(na500_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a504_5 ( .OUT(na504_2), .CLK(na367_1), .EN(na14_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na504_2_i) );
// C_AND/D//AND/D      x103y11     80'h00_EA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a532_1 ( .OUT(na532_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na370_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a532_2 ( .OUT(na532_1), .CLK(na367_1), .EN(na97_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na532_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a532_4 ( .OUT(na532_2_i), .IN1(1'b1), .IN2(na370_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a532_5 ( .OUT(na532_2), .CLK(na367_1), .EN(na97_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na532_2_i) );
// C_AND/D//AND/D      x105y16     80'h00_EA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a533_1 ( .OUT(na533_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na375_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a533_2 ( .OUT(na533_1), .CLK(na367_1), .EN(na97_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na533_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a533_4 ( .OUT(na533_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na375_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a533_5 ( .OUT(na533_2), .CLK(na367_1), .EN(na97_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na533_2_i) );
// C_AND/D//AND/D      x110y27     80'h00_EA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a534_1 ( .OUT(na534_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na376_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a534_2 ( .OUT(na534_1), .CLK(na367_1), .EN(na97_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na534_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a534_4 ( .OUT(na534_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na376_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a534_5 ( .OUT(na534_2), .CLK(na367_1), .EN(na97_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na534_2_i) );
// C_AND/D//AND/D      x105y27     80'h00_EA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a538_1 ( .OUT(na538_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na374_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a538_2 ( .OUT(na538_1), .CLK(na367_1), .EN(na97_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na538_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a538_4 ( .OUT(na538_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na374_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a538_5 ( .OUT(na538_2), .CLK(na367_1), .EN(na97_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na538_2_i) );
// C_AND/D///      x90y30     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a539_1 ( .OUT(na539_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na82_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a539_2 ( .OUT(na539_1), .CLK(na367_1), .EN(na283_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na539_1_i) );
// C_///AND/D      x89y26     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a540_4 ( .OUT(na540_2_i), .IN1(1'b1), .IN2(na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a540_5 ( .OUT(na540_2), .CLK(na367_1), .EN(na285_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na540_2_i) );
// C_AND/D//AND/D      x93y29     80'h00_EA00_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a542_1 ( .OUT(na542_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na225_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a542_2 ( .OUT(na542_1), .CLK(na367_1), .EN(na46_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na542_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a542_4 ( .OUT(na542_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na550_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a542_5 ( .OUT(na542_2), .CLK(na367_1), .EN(na46_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na542_2_i) );
// C_///AND/D      x95y21     80'h00_EA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a543_4 ( .OUT(na543_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na550_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a543_5 ( .OUT(na543_2), .CLK(na367_1), .EN(na46_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na543_2_i) );
// C_AND/D//AND/D      x95y28     80'h00_EA00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a546_1 ( .OUT(na546_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na548_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a546_2 ( .OUT(na546_1), .CLK(na367_1), .EN(na46_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na546_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a546_4 ( .OUT(na546_2_i), .IN1(na542_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a546_5 ( .OUT(na546_2), .CLK(na367_1), .EN(na46_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na546_2_i) );
// C_///AND/D      x96y27     80'h00_EA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a547_4 ( .OUT(na547_2_i), .IN1(na542_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a547_5 ( .OUT(na547_2), .CLK(na367_1), .EN(na46_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na547_2_i) );
// C_AND/D///      x93y26     80'h00_EA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a548_1 ( .OUT(na548_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na546_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a548_2 ( .OUT(na548_1), .CLK(na367_1), .EN(na46_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na548_1_i) );
// C_AND/D//AND/D      x96y26     80'h00_EA00_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a550_1 ( .OUT(na550_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na546_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a550_2 ( .OUT(na550_1), .CLK(na367_1), .EN(na46_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na550_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a550_4 ( .OUT(na550_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na547_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a550_5 ( .OUT(na550_2), .CLK(na367_1), .EN(na46_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na550_2_i) );
// C_///AND/D      x91y27     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a556_4 ( .OUT(na556_2_i), .IN1(1'b1), .IN2(na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a556_5 ( .OUT(na556_2), .CLK(na367_1), .EN(na286_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na556_2_i) );
// C_AND/D//AND/D      x107y30     80'h00_EA00_80_0000_0C88_CFF3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a567_1 ( .OUT(na567_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na348_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a567_2 ( .OUT(na567_1), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na567_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a567_4 ( .OUT(na567_2_i), .IN1(1'b1), .IN2(~na567_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a567_5 ( .OUT(na567_2), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na567_2_i) );
// C_AND/D///      x107y31     80'h00_EA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a569_1 ( .OUT(na569_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na350_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a569_2 ( .OUT(na569_1), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na569_1_i) );
// C_///AND/D      x107y25     80'h00_EA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a573_4 ( .OUT(na573_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na354_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a573_5 ( .OUT(na573_2), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na573_2_i) );
// C_///AND/D      x110y29     80'h00_EA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a575_4 ( .OUT(na575_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na356_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a575_5 ( .OUT(na575_2), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na575_2_i) );
// C_AND/D//AND/D      x109y32     80'h00_EA00_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a577_1 ( .OUT(na577_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na344_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a577_2 ( .OUT(na577_1), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na577_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a577_4 ( .OUT(na577_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na352_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a577_5 ( .OUT(na577_2), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na577_2_i) );
// C_///AND/D      x107y31     80'h00_EA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a579_4 ( .OUT(na579_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na346_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a579_5 ( .OUT(na579_2), .CLK(na367_1), .EN(na272_2), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na579_2_i) );
// C_AND/D///      x95y30     80'h00_E600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a581_1 ( .OUT(na581_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na604_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a581_2 ( .OUT(na581_1), .CLK(na367_1), .EN(~na139_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na581_1_i) );
// C_///AND/D      x96y32     80'h00_E600_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a582_4 ( .OUT(na582_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na605_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a582_5 ( .OUT(na582_2), .CLK(na367_1), .EN(~na139_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na582_2_i) );
// C_AND/D///      x100y31     80'h00_E600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a583_1 ( .OUT(na583_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na606_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a583_2 ( .OUT(na583_1), .CLK(na367_1), .EN(~na139_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na583_1_i) );
// C_AND/D///      x99y27     80'h00_E600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a584_1 ( .OUT(na584_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na607_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a584_2 ( .OUT(na584_1), .CLK(na367_1), .EN(~na139_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na584_1_i) );
// C_AND/D///      x97y30     80'h00_E600_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a585_1 ( .OUT(na585_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na608_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a585_2 ( .OUT(na585_1), .CLK(na367_1), .EN(~na139_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na585_1_i) );
// C_///AND/D      x100y31     80'h00_E600_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a586_4 ( .OUT(na586_2_i), .IN1(1'b1), .IN2(na609_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a586_5 ( .OUT(na586_2), .CLK(na367_1), .EN(~na139_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na586_2_i) );
// C_AND/D///      x98y28     80'h00_E600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a587_1 ( .OUT(na587_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na610_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a587_2 ( .OUT(na587_1), .CLK(na367_1), .EN(~na139_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na587_1_i) );
// C_///AND/D      x96y22     80'h00_E600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a588_4 ( .OUT(na588_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na611_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a588_5 ( .OUT(na588_2), .CLK(na367_1), .EN(~na139_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na588_2_i) );
// C_AND/DST///      x109y8     80'h20_BA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a590_1 ( .OUT(na590_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na266_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'b1_0100_0000)) 
           _a590_2 ( .OUT(na590_1), .CLK(na367_1), .EN(na267_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na590_1_i) );
// C_AND/D///      x95y27     80'h00_EA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a591_1 ( .OUT(na591_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na604_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a591_2 ( .OUT(na591_1), .CLK(na367_1), .EN(na128_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na591_1_i) );
// C_AND/D///      x95y31     80'h00_EA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a592_1 ( .OUT(na592_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na605_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a592_2 ( .OUT(na592_1), .CLK(na367_1), .EN(na128_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na592_1_i) );
// C_///AND/D      x98y29     80'h00_EA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a593_4 ( .OUT(na593_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na606_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a593_5 ( .OUT(na593_2), .CLK(na367_1), .EN(na128_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na593_2_i) );
// C_AND/D///      x100y29     80'h00_EA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a594_1 ( .OUT(na594_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na607_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a594_2 ( .OUT(na594_1), .CLK(na367_1), .EN(na128_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na594_1_i) );
// C_///AND/D      x101y31     80'h00_EA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a595_4 ( .OUT(na595_2_i), .IN1(1'b1), .IN2(na608_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a595_5 ( .OUT(na595_2), .CLK(na367_1), .EN(na128_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na595_2_i) );
// C_///AND/D      x95y29     80'h00_EA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a596_4 ( .OUT(na596_2_i), .IN1(1'b1), .IN2(na609_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a596_5 ( .OUT(na596_2), .CLK(na367_1), .EN(na128_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na596_2_i) );
// C_///AND/D      x100y29     80'h00_EA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a597_4 ( .OUT(na597_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na610_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a597_5 ( .OUT(na597_2), .CLK(na367_1), .EN(na128_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na597_2_i) );
// C_AND/D///      x100y26     80'h00_EA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a598_1 ( .OUT(na598_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na611_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a598_2 ( .OUT(na598_1), .CLK(na367_1), .EN(na128_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na598_1_i) );
// C_MX4b////      x88y30     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a600_1 ( .OUT(na600_1), .IN1(1'b1), .IN2(na843_2), .IN3(1'b1), .IN4(~na409_2), .IN5(na556_2), .IN6(na540_2), .IN7(na368_2),
                     .IN8(na366_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x90y31     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a601_1 ( .OUT(na601_1), .IN1(1'b1), .IN2(~na843_2), .IN3(1'b1), .IN4(~na409_2), .IN5(na494_2), .IN6(na492_2), .IN7(na493_1),
                     .IN8(na539_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000050)) 
           _a602 ( .Y(na602_1), .I(arst_n) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a603 ( .Y(na603_1), .I(clk) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a604 ( .Y(na604_1), .O(io_psram_data0), .A(na766_10), .EN(na767_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a605 ( .Y(na605_1), .O(io_psram_data1), .A(na768_10), .EN(na769_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a606 ( .Y(na606_1), .O(io_psram_data2), .A(na770_10), .EN(na771_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a607 ( .Y(na607_1), .O(io_psram_data3), .A(na772_10), .EN(na773_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a608 ( .Y(na608_1), .O(io_psram_data4), .A(na774_10), .EN(na775_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a609 ( .Y(na609_1), .O(io_psram_data5), .A(na776_10), .EN(na777_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a610 ( .Y(na610_1), .O(io_psram_data6), .A(na778_10), .EN(na779_10) );
CPE_IOBF   #(.BUF_CFG (72'h000001000100060910)) 
           _a611 ( .Y(na611_1), .O(io_psram_data7), .A(na780_10), .EN(na781_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a612 ( .O(led), .A(na782_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a613 ( .O(o_psram_csn), .A(na783_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a614 ( .O(o_psram_sclk), .A(na784_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a615 ( .O(sent), .A(na785_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a616 ( .O(tick_1us), .A(na786_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a617 ( .Y(na617_1), .I(uart_rx) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a618 ( .O(uart_tx), .A(na787_10) );
// C_AND////      x103y27     80'h00_0018_00_0000_0888_1223
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a619_1 ( .OUT(na619_1), .IN1(1'b1), .IN2(~na442_1), .IN3(na234_1), .IN4(~na280_2), .IN5(na4_1), .IN6(~na442_2), .IN7(~na443_1),
                     .IN8(~na444_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/DST      x91y10     80'h20_BA00_80_0000_0C08_FF00
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a620_4 ( .OUT(na620_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_DST      #(.CPE_CFG (9'b1_0100_0100)) 
           _a620_5 ( .OUT(na620_2), .CLK(na367_1), .EN(na277_1), .SR(na602_1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na620_2_i) );
// C_/C_0_1///      x98y9     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a621_2 ( .OUT(na621_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a621_6 ( .COUTY1(na621_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na621_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x97y11     80'h00_0018_00_0000_0CEE_EC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a622_1 ( .OUT(na622_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na500_1), .IN7(na221_2), .IN8(na503_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x95y9     80'h00_0018_00_0000_0888_5341
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a624_1 ( .OUT(na624_1), .IN1(~na504_2), .IN2(~na501_1), .IN3(~na502_1), .IN4(na20_1), .IN5(1'b1), .IN6(~na501_2), .IN7(~na502_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x99y11     80'h00_0018_00_0000_0888_F53B
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a625_1 ( .OUT(na625_1), .IN1(na849_2), .IN2(~na237_1), .IN3(1'b0), .IN4(~na25_1), .IN5(~na21_2), .IN6(1'b0), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x95y13     80'h00_0018_00_0000_0888_F5B5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a629_1 ( .OUT(na629_1), .IN1(~na42_1), .IN2(1'b0), .IN3(na799_2), .IN4(~na631_1), .IN5(~na42_2), .IN6(1'b0), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x94y15     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a630_4 ( .OUT(na630_2), .IN1(~na543_2), .IN2(1'b1), .IN3(1'b1), .IN4(na752_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x92y10     80'h00_0018_00_0000_0CEE_A300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a631_1 ( .OUT(na631_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na31_2), .IN7(na630_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x94y17     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a633_1 ( .OUT(na633_1), .IN1(~na45_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na837_2), .IN6(na46_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x94y12     80'h00_0018_00_0000_0888_F373
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a634_1 ( .OUT(na634_1), .IN1(1'b0), .IN2(~na49_1), .IN3(~na53_2), .IN4(~na631_1), .IN5(1'b0), .IN6(~na49_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x91y12     80'h00_0018_00_0000_0888_7F53
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a639_1 ( .OUT(na639_1), .IN1(1'b0), .IN2(~na49_1), .IN3(~na55_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(~na53_1), .IN8(~na631_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x95y16     80'h00_0018_00_0000_0888_5FB3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a644_1 ( .OUT(na644_1), .IN1(1'b0), .IN2(~na49_1), .IN3(na801_2), .IN4(~na631_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na58_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y27     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a650_4 ( .OUT(na650_2), .IN1(na66_2), .IN2(na93_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x92y30     80'h00_0078_00_0000_0C88_AAAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a651_1 ( .OUT(na651_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na10_2), .IN6(1'b1), .IN7(na8_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a651_4 ( .OUT(na651_2), .IN1(1'b1), .IN2(na546_2), .IN3(na103_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x93y20     80'h00_0018_00_0000_0EEE_EA5D
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a652_1 ( .OUT(na652_1), .IN1(~na98_1), .IN2(na41_2), .IN3(~na225_1), .IN4(1'b0), .IN5(na56_1), .IN6(1'b0), .IN7(na53_1),
                     .IN8(na800_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x93y32     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a655_1 ( .OUT(na655_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na100_1), .IN6(1'b1), .IN7(na547_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x89y27     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a656_4 ( .OUT(na656_2), .IN1(~na104_1), .IN2(~na548_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x94y20     80'h00_0018_00_0000_0CEE_7300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a660_1 ( .OUT(na660_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na90_2), .IN7(~na805_2), .IN8(~na89_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x98y21     80'h00_0018_00_0000_0888_2435
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a667_1 ( .OUT(na667_1), .IN1(~na125_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na155_1), .IN5(~na127_1), .IN6(na157_1), .IN7(na156_2),
                     .IN8(~na133_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x99y26     80'h00_0018_00_0000_0C66_3C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a671_1 ( .OUT(na671_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na295_1), .IN7(1'b0), .IN8(~na108_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x98y19     80'h00_0018_00_0040_0A64_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a679_1 ( .OUT(na679_1), .IN1(1'b1), .IN2(~na153_2), .IN3(1'b1), .IN4(na825_2), .IN5(1'b0), .IN6(na832_2), .IN7(~na161_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x99y22     80'h00_0060_00_0000_0C08_FF52
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a680_4 ( .OUT(na680_2), .IN1(na137_2), .IN2(~na150_2), .IN3(~na63_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y17     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a681_4 ( .OUT(na681_2), .IN1(1'b1), .IN2(1'b1), .IN3(na62_2), .IN4(~na164_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x101y21     80'h00_0078_00_0000_0C88_75AE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a683_1 ( .OUT(na683_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na130_2), .IN6(1'b0), .IN7(~na812_2), .IN8(~na111_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a683_4 ( .OUT(na683_2), .IN1(na130_1), .IN2(na114_1), .IN3(na62_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x105y12     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a685_1 ( .OUT(na685_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na446_2), .IN6(1'b0), .IN7(~na173_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x106y15     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a686_1 ( .OUT(na686_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na466_1), .IN6(~na186_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x105y15     80'h00_0060_00_0000_0C0E_FF70
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a694_4 ( .OUT(na694_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na474_2), .IN4(~na817_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x107y15     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a695_1 ( .OUT(na695_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na168_1), .IN8(na488_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y11     80'h00_0018_00_0000_0888_F541
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a696_1 ( .OUT(na696_1), .IN1(~na698_1), .IN2(~na188_1), .IN3(~na187_2), .IN4(na697_1), .IN5(~na698_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x102y14     80'h00_0018_00_0000_0CEE_B000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a697_1 ( .OUT(na697_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na173_2), .IN8(~na455_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x103y13     80'h00_0078_00_0000_0C88_C3C3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a698_1 ( .OUT(na698_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na186_2), .IN7(1'b1), .IN8(na463_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a698_4 ( .OUT(na698_2), .IN1(1'b1), .IN2(~na186_1), .IN3(1'b1), .IN4(na463_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x108y14     80'h00_0060_00_0000_0C0E_FF53
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a702_4 ( .OUT(na702_2), .IN1(1'b0), .IN2(~na475_1), .IN3(~na121_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x108y11     80'h00_0078_00_0000_0C88_AA8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a703_1 ( .OUT(na703_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na489_1), .IN6(1'b1), .IN7(na168_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a703_4 ( .OUT(na703_2), .IN1(1'b1), .IN2(1'b1), .IN3(na459_1), .IN4(na190_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x104y17     80'h00_0018_00_0000_0888_1C14
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a704_1 ( .OUT(na704_1), .IN1(~na821_2), .IN2(na705_1), .IN3(~na123_2), .IN4(~na706_2), .IN5(1'b1), .IN6(na705_2), .IN7(~na823_2),
                     .IN8(~na706_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x107y20     80'h00_0078_00_0000_0CEE_0D35
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a705_1 ( .OUT(na705_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na464_1), .IN6(na186_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a705_4 ( .OUT(na705_2), .IN1(~na683_2), .IN2(1'b0), .IN3(1'b0), .IN4(~na452_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x106y18     80'h00_0078_00_0000_0C88_4FAA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a706_1 ( .OUT(na706_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na173_2), .IN8(na456_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a706_4 ( .OUT(na706_2), .IN1(na448_2), .IN2(1'b1), .IN3(na173_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x109y15     80'h00_0078_00_0000_0CEE_3C70
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a710_1 ( .OUT(na710_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na186_2), .IN7(1'b0), .IN8(~na468_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a710_4 ( .OUT(na710_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na121_1), .IN4(~na476_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x110y14     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a711_4 ( .OUT(na711_2), .IN1(na460_2), .IN2(1'b1), .IN3(1'b1), .IN4(na190_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x108y12     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a713_4 ( .OUT(na713_2), .IN1(1'b1), .IN2(na490_1), .IN3(na168_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x105y24     80'h00_0018_00_0000_0888_3352
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a714_1 ( .OUT(na714_1), .IN1(na715_1), .IN2(~na716_1), .IN3(~na202_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na716_2), .IN7(1'b1),
                     .IN8(~na203_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x105y23     80'h00_0018_00_0000_0CEE_B000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a715_1 ( .OUT(na715_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na173_2), .IN8(~na457_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x103y24     80'h00_0078_00_0000_0C88_F2F2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a716_1 ( .OUT(na716_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na465_2), .IN6(~na186_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a716_4 ( .OUT(na716_2), .IN1(na465_1), .IN2(~na186_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x111y19     80'h00_0060_00_0000_0C0E_FF53
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a718_4 ( .OUT(na718_2), .IN1(1'b0), .IN2(~na477_1), .IN3(~na121_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x109y17     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a719_1 ( .OUT(na719_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na491_1), .IN7(na168_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x106y11     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a720_4 ( .OUT(na720_2), .IN1(~na470_2), .IN2(1'b0), .IN3(~na121_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x107y11     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a721_1 ( .OUT(na721_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na168_1), .IN8(na484_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x106y10     80'h00_0018_00_0000_0CEE_5500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a723_1 ( .OUT(na723_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na471_1), .IN6(1'b0), .IN7(~na121_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x108y9     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a724_4 ( .OUT(na724_2), .IN1(na485_2), .IN2(1'b1), .IN3(na168_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x110y13     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a726_1 ( .OUT(na726_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na472_2), .IN7(~na121_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x110y14     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a727_1 ( .OUT(na727_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na486_2), .IN6(1'b1), .IN7(na168_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x107y17     80'h00_0060_00_0000_0C0E_FF55
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a729_4 ( .OUT(na729_2), .IN1(~na473_2), .IN2(1'b0), .IN3(~na121_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x109y17     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a730_4 ( .OUT(na730_2), .IN1(1'b1), .IN2(na834_2), .IN3(na487_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x98y13     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a736_4 ( .OUT(na736_2), .IN1(na140_1), .IN2(na295_1), .IN3(na62_1), .IN4(na108_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x97y14     80'h00_0078_00_0000_0C88_F441
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a737_1 ( .OUT(na737_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na167_1), .IN6(na150_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a737_4 ( .OUT(na737_2), .IN1(~na141_1), .IN2(~na295_1), .IN3(~na161_1), .IN4(na108_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x104y19     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a746_4 ( .OUT(na746_2), .IN1(na97_2), .IN2(~na258_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x94y24     80'h00_0078_00_0000_0C88_332A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a752_1 ( .OUT(na752_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na548_1), .IN7(1'b1), .IN8(~na550_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a752_4 ( .OUT(na752_2), .IN1(na10_2), .IN2(1'b1), .IN3(na8_1), .IN4(~na550_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x107y9     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a753_1 ( .OUT(na753_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na262_2), .IN6(1'b1), .IN7(1'b1), .IN8(na266_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y26     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a755_1 ( .OUT(na755_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na150_2), .IN7(na62_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x106y31     80'h00_0018_00_0000_0EEE_3375
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a757_1 ( .OUT(na757_1), .IN1(~na579_2), .IN2(1'b0), .IN3(~na575_2), .IN4(~na356_1), .IN5(1'b0), .IN6(~na567_2), .IN7(1'b0),
                     .IN8(~na758_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x108y32     80'h00_0018_00_0000_0888_2112
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a758_1 ( .OUT(na758_1), .IN1(na276_1), .IN2(~na577_1), .IN3(~na845_2), .IN4(~na352_1), .IN5(~na573_2), .IN6(~na577_2), .IN7(na344_1),
                     .IN8(~na846_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x101y13     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a759_4 ( .OUT(na759_2), .IN1(~na262_2), .IN2(~na226_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x99y19     80'h00_0018_00_0000_0C88_EAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a762_1 ( .OUT(na762_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na293_1), .IN6(1'b0), .IN7(na62_1), .IN8(na111_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x101y19     80'h00_0018_00_0000_0888_2412
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a765_1 ( .OUT(na765_1), .IN1(na296_2), .IN2(~na118_2), .IN3(~na173_1), .IN4(~na147_2), .IN5(~na683_2), .IN6(na157_1), .IN7(na156_2),
                     .IN8(~na190_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x121y1     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a766_4 ( .OUT(na766_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na208_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a766_6 ( .RAM_O2(na766_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na766_2), .COMP_OUT(1'b0) );
// C_///AND/      x122y1     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a767_4 ( .OUT(na767_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na266_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a767_6 ( .RAM_O2(na767_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na767_2), .COMP_OUT(1'b0) );
// C_///AND/      x123y1     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a768_4 ( .OUT(na768_2), .IN1(na210_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a768_6 ( .RAM_O2(na768_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na768_2), .COMP_OUT(1'b0) );
// C_///AND/      x124y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a769_4 ( .OUT(na769_2), .IN1(1'b1), .IN2(na590_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a769_6 ( .RAM_O2(na769_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na769_2), .COMP_OUT(1'b0) );
// C_///AND/      x125y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a770_4 ( .OUT(na770_2), .IN1(1'b1), .IN2(na212_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a770_6 ( .RAM_O2(na770_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na770_2), .COMP_OUT(1'b0) );
// C_///AND/      x126y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a771_4 ( .OUT(na771_2), .IN1(1'b1), .IN2(na590_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a771_6 ( .RAM_O2(na771_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na771_2), .COMP_OUT(1'b0) );
// C_///AND/      x127y1     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a772_4 ( .OUT(na772_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na214_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a772_6 ( .RAM_O2(na772_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na772_2), .COMP_OUT(1'b0) );
// C_///AND/      x128y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a773_4 ( .OUT(na773_2), .IN1(1'b1), .IN2(na590_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a773_6 ( .RAM_O2(na773_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na773_2), .COMP_OUT(1'b0) );
// C_///AND/      x129y1     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a774_4 ( .OUT(na774_2), .IN1(na169_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a774_6 ( .RAM_O2(na774_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na774_2), .COMP_OUT(1'b0) );
// C_///AND/      x130y1     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a775_4 ( .OUT(na775_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na266_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a775_6 ( .RAM_O2(na775_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na775_2), .COMP_OUT(1'b0) );
// C_///AND/      x131y1     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a776_4 ( .OUT(na776_2), .IN1(na182_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a776_6 ( .RAM_O2(na776_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na776_2), .COMP_OUT(1'b0) );
// C_///AND/      x132y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a777_4 ( .OUT(na777_2), .IN1(1'b1), .IN2(na590_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a777_6 ( .RAM_O2(na777_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na777_2), .COMP_OUT(1'b0) );
// C_///AND/      x133y1     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a778_4 ( .OUT(na778_2), .IN1(1'b1), .IN2(1'b1), .IN3(na192_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a778_6 ( .RAM_O2(na778_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na778_2), .COMP_OUT(1'b0) );
// C_///AND/      x134y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a779_4 ( .OUT(na779_2), .IN1(1'b1), .IN2(na590_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a779_6 ( .RAM_O2(na779_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na779_2), .COMP_OUT(1'b0) );
// C_///AND/      x135y1     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a780_4 ( .OUT(na780_2), .IN1(1'b1), .IN2(1'b1), .IN3(na199_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a780_6 ( .RAM_O2(na780_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na780_2), .COMP_OUT(1'b0) );
// C_///AND/      x136y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a781_4 ( .OUT(na781_2), .IN1(1'b1), .IN2(na590_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a781_6 ( .RAM_O2(na781_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na781_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y95     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a782_4 ( .OUT(na782_2), .IN1(na96_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a782_6 ( .RAM_O2(na782_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na782_2), .COMP_OUT(1'b0) );
// C_///AND/      x117y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a783_4 ( .OUT(na783_2), .IN1(1'b1), .IN2(na226_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a783_6 ( .RAM_O2(na783_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na783_2), .COMP_OUT(1'b0) );
// C_///AND/      x119y1     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a784_4 ( .OUT(na784_2), .IN1(1'b1), .IN2(na106_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a784_6 ( .RAM_O2(na784_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na784_2), .COMP_OUT(1'b0) );
// C_///AND/      x160y73     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a785_4 ( .OUT(na785_2), .IN1(1'b1), .IN2(na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a785_6 ( .RAM_O2(na785_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na785_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y45     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a786_4 ( .OUT(na786_2), .IN1(1'b1), .IN2(na31_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a786_6 ( .RAM_O2(na786_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na786_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y51     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a787_4 ( .OUT(na787_2), .IN1(1'b1), .IN2(na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a787_6 ( .RAM_O2(na787_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                     .OUT2(na787_2), .COMP_OUT(1'b0) );
// C_////Bridge      x101y28     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a788_5 ( .OUT(na788_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na6_1) );
// C_////Bridge      x98y7     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a789_5 ( .OUT(na789_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na11_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y8     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a790_5 ( .OUT(na790_2), .IN1(na21_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y7     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a791_5 ( .OUT(na791_2), .IN1(1'b0), .IN2(1'b0), .IN3(na26_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x92y12     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a792_5 ( .OUT(na792_2), .IN1(1'b0), .IN2(na31_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y16     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a793_5 ( .OUT(na793_2), .IN1(1'b0), .IN2(na31_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y9     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a794_5 ( .OUT(na794_2), .IN1(1'b0), .IN2(1'b0), .IN3(na33_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y25     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a795_5 ( .OUT(na795_2), .IN1(1'b0), .IN2(na38_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y19     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a796_5 ( .OUT(na796_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na39_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y25     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a797_5 ( .OUT(na797_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na39_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y23     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a798_5 ( .OUT(na798_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na39_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y11     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a799_5 ( .OUT(na799_2), .IN1(1'b0), .IN2(na41_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y18     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a800_5 ( .OUT(na800_2), .IN1(1'b0), .IN2(1'b0), .IN3(na53_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x96y13     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a801_5 ( .OUT(na801_2), .IN1(na56_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y6     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a802_5 ( .OUT(na802_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na61_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y19     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a803_5 ( .OUT(na803_2), .IN1(1'b0), .IN2(1'b0), .IN3(na62_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y30     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a804_5 ( .OUT(na804_2), .IN1(1'b0), .IN2(1'b0), .IN3(na64_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x88y17     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a805_5 ( .OUT(na805_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na89_2) );
// C_////Bridge      x104y21     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a806_5 ( .OUT(na806_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na108_1) );
// C_////Bridge      x102y19     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a807_5 ( .OUT(na807_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na110_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y18     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a808_5 ( .OUT(na808_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na111_2) );
// C_////Bridge      x102y16     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a809_5 ( .OUT(na809_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na112_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y15     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a810_5 ( .OUT(na810_2), .IN1(1'b0), .IN2(na114_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y13     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a811_5 ( .OUT(na811_2), .IN1(1'b0), .IN2(na114_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x106y19     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a812_5 ( .OUT(na812_2), .IN1(1'b0), .IN2(na114_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y15     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a813_5 ( .OUT(na813_2), .IN1(na117_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y19     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a814_5 ( .OUT(na814_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na119_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x105y18     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a815_5 ( .OUT(na815_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na119_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y19     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a816_5 ( .OUT(na816_2), .IN1(1'b0), .IN2(1'b0), .IN3(na120_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y14     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a817_5 ( .OUT(na817_2), .IN1(1'b0), .IN2(1'b0), .IN3(na121_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y21     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a818_5 ( .OUT(na818_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na123_2), .IN8(1'b0) );
// C_////Bridge      x104y15     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a819_5 ( .OUT(na819_2), .IN1(na130_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y14     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a820_5 ( .OUT(na820_2), .IN1(na130_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x107y15     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a821_5 ( .OUT(na821_2), .IN1(1'b0), .IN2(na136_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y15     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a822_5 ( .OUT(na822_2), .IN1(1'b0), .IN2(na136_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x108y17     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a823_5 ( .OUT(na823_2), .IN1(1'b0), .IN2(na136_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y16     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a824_5 ( .OUT(na824_2), .IN1(na141_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x100y20     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a825_5 ( .OUT(na825_2), .IN1(na141_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x102y11     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a826_5 ( .OUT(na826_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na144_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y14     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a827_5 ( .OUT(na827_2), .IN1(na146_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x101y20     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a828_5 ( .OUT(na828_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na147_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x98y15     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a829_5 ( .OUT(na829_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na148_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y24     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a830_5 ( .OUT(na830_2), .IN1(1'b0), .IN2(na150_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y21     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a831_5 ( .OUT(na831_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na155_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y18     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a832_5 ( .OUT(na832_2), .IN1(1'b0), .IN2(1'b0), .IN3(na161_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x104y16     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a833_5 ( .OUT(na833_2), .IN1(1'b0), .IN2(1'b0), .IN3(na161_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x111y18     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a834_5 ( .OUT(na834_2), .IN1(1'b0), .IN2(1'b0), .IN3(na168_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x90y21     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a835_5 ( .OUT(na835_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na216_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y23     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a836_5 ( .OUT(na836_2), .IN1(1'b0), .IN2(1'b0), .IN3(na225_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x95y15     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a837_5 ( .OUT(na837_2), .IN1(1'b0), .IN2(1'b0), .IN3(na235_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x112y22     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a838_5 ( .OUT(na838_2), .IN1(1'b0), .IN2(na238_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y21     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a839_5 ( .OUT(na839_2), .IN1(na240_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x109y5     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a840_5 ( .OUT(na840_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na266_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y13     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a841_5 ( .OUT(na841_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na280_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y21     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a842_5 ( .OUT(na842_2), .IN1(1'b0), .IN2(1'b0), .IN3(na288_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x91y30     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a843_5 ( .OUT(na843_2), .IN1(1'b0), .IN2(1'b0), .IN3(na318_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x89y30     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a844_5 ( .OUT(na844_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na320_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y31     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a845_5 ( .OUT(na845_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na346_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x110y32     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a846_5 ( .OUT(na846_2), .IN1(1'b0), .IN2(1'b0), .IN3(na354_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x93y26     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a847_5 ( .OUT(na847_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na409_2) );
// C_////Bridge      x109y24     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a848_5 ( .OUT(na848_2), .IN1(na438_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x99y9     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a849_5 ( .OUT(na849_2), .IN1(1'b0), .IN2(1'b0), .IN3(na497_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x100y15     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a850_5 ( .OUT(na850_2), .IN1(na683_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x103y17     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a851_5 ( .OUT(na851_2), .IN1(1'b0), .IN2(na737_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x97y19     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a852_5 ( .OUT(na852_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na752_1) );
endmodule
