//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 January 2025)
//  Compile Time: 2025-03-05 10:25:39
//  Program Run:  2025-03-05 13:06:38
//  Program Call: /home/tarik/Downloads/cc-toolchain-linux/bin/p_r/p_r -A 1 -i corescore_0_synth.v -o corescore_0 -lib ccag -cCP --verbose -tm 1 -ccf src/corescore_0/data/cc_gatemate.ccf 
//  File Type:    Verilog

// Gatecount:   2880
module corescore_0 (i_clk , i_rstn ,
       o_uart_tx 
       ) ;

input  i_clk;
input  i_rstn;

output o_uart_tx;



wire i_clk;
wire na2_1;
wire na2_2;
wire na3_1;
wire na4_1;
wire na7_2;
wire na8_1;
wire na9_1;
wire na9_2;
wire i_rstn;
wire na11_1;
wire na12_1;
wire na15_2;
wire na16_1;
wire na17_1;
wire na17_2;
wire na19_1;
wire na21_1;
wire na22_1;
wire na22_2;
wire na24_1;
wire na25_2;
wire na26_1;
wire na27_1;
wire na27_2;
wire na28_1;
wire na30_1;
wire na30_1_i;
wire na31_2;
wire na32_1;
wire na32_1_i;
wire na33_1;
wire na34_1;
wire na34_1_i;
wire na35_1;
wire na35_1_i;
wire na36_1;
wire na36_1_i;
wire na37_1;
wire na37_1_i;
wire na38_1;
wire na38_1_i;
wire na38_2;
wire na38_2_i;
wire na39_1;
wire na39_1_i;
wire na40_1;
wire na40_1_i;
wire na41_1;
wire na41_1_i;
wire na42_1;
wire na42_1_i;
wire na43_1;
wire na43_1_i;
wire na44_1;
wire na44_1_i;
wire na45_1;
wire na45_1_i;
wire na46_1;
wire na46_1_i;
wire na47_1;
wire na47_1_i;
wire na48_1;
wire na48_1_i;
wire na49_1;
wire na49_1_i;
wire na50_1;
wire na50_1_i;
wire na51_1;
wire na51_1_i;
wire na52_1;
wire na52_1_i;
wire na53_1;
wire na53_1_i;
wire na54_2;
wire na55_1;
wire na55_2;
wire na56_1;
wire na56_1_i;
wire na57_1;
wire na57_1_i;
wire na58_1;
wire na58_1_i;
wire na59_1;
wire na59_1_i;
wire na60_1;
wire na60_1_i;
wire na61_1;
wire na61_1_i;
wire na62_1;
wire na62_1_i;
wire na63_1;
wire na63_1_i;
wire na64_1;
wire na64_1_i;
wire na65_1;
wire na65_1_i;
wire na66_1;
wire na66_1_i;
wire na67_1;
wire na67_1_i;
wire na68_1;
wire na68_1_i;
wire na69_1;
wire na69_1_i;
wire na70_1;
wire na70_1_i;
wire na71_1;
wire na71_1_i;
wire na72_1;
wire na72_1_i;
wire na73_1;
wire na73_1_i;
wire na75_1;
wire na75_1_i;
wire na76_1;
wire na76_1_i;
wire na76_2;
wire na76_2_i;
wire na78_1;
wire na78_1_i;
wire na78_2;
wire na78_2_i;
wire na79_1;
wire na79_1_i;
wire na79_2;
wire na79_2_i;
wire na80_1;
wire na80_1_i;
wire na81_1;
wire na83_2;
wire na84_2;
wire na84_2_i;
wire na85_1;
wire na85_1_i;
wire na85_2;
wire na85_2_i;
wire na87_1;
wire na87_1_i;
wire na88_1;
wire na88_1_i;
wire na88_2;
wire na88_2_i;
wire na89_1;
wire na89_1_i;
wire na89_2;
wire na89_2_i;
wire na90_1;
wire na90_2;
wire na91_1;
wire na92_1;
wire na93_1;
wire na94_1;
wire na94_2;
wire na95_1;
wire na95_2;
wire na98_1;
wire na103_1;
wire na103_1_i;
wire na104_1;
wire na104_1_i;
wire na105_1;
wire na105_1_i;
wire na107_1;
wire na107_1_i;
wire na108_1;
wire na108_1_i;
wire na109_1;
wire na109_1_i;
wire na110_1;
wire na110_1_i;
wire na111_1;
wire na111_1_i;
wire na112_1;
wire na112_1_i;
wire na113_1;
wire na113_1_i;
wire na114_1;
wire na114_1_i;
wire na115_1;
wire na115_1_i;
wire na117_1;
wire na117_2;
wire na118_1;
wire na118_1_i;
wire na119_1;
wire na119_1_i;
wire na120_2;
wire na121_2;
wire na122_1;
wire na122_2;
wire na123_1;
wire na123_1_i;
wire na124_1;
wire na124_1_i;
wire na125_1;
wire na125_1_i;
wire na126_1;
wire na126_1_i;
wire na127_1;
wire na127_1_i;
wire na128_1;
wire na128_1_i;
wire na129_1;
wire na129_1_i;
wire na130_1;
wire na130_1_i;
wire na131_1;
wire na131_1_i;
wire na132_1;
wire na132_1_i;
wire na133_1;
wire na133_1_i;
wire na134_1;
wire na134_1_i;
wire na135_1;
wire na135_1_i;
wire na136_1;
wire na136_1_i;
wire na137_2;
wire na138_1;
wire na139_1;
wire na143_1;
wire na145_1;
wire na146_1;
wire na153_1;
wire na153_1_i;
wire na154_1;
wire na154_1_i;
wire na155_2;
wire na156_1;
wire na157_1;
wire na157_1_i;
wire na158_1;
wire na158_1_i;
wire na159_1;
wire na159_1_i;
wire na160_1;
wire na160_1_i;
wire na161_1;
wire na161_1_i;
wire na162_1;
wire na162_1_i;
wire na163_1;
wire na163_1_i;
wire na164_1;
wire na164_1_i;
wire na165_1;
wire na165_1_i;
wire na166_1;
wire na166_1_i;
wire na167_1;
wire na167_1_i;
wire na168_1;
wire na168_1_i;
wire na169_1;
wire na169_1_i;
wire na170_1;
wire na170_1_i;
wire na171_1;
wire na171_1_i;
wire na173_1;
wire na173_1_i;
wire na174_1;
wire na174_1_i;
wire na175_1;
wire na176_2;
wire na178_1;
wire na179_1;
wire na180_1;
wire na181_1;
wire na182_1;
wire na187_2;
wire na188_1;
wire na189_2;
wire na190_1;
wire na190_1_i;
wire na190_2;
wire na190_2_i;
wire na192_1;
wire na192_1_i;
wire na192_2;
wire na192_2_i;
wire na193_1;
wire na193_1_i;
wire na193_2;
wire na193_2_i;
wire na194_1;
wire na196_2;
wire na197_1;
wire na197_1_i;
wire na198_1;
wire na198_2;
wire na200_1;
wire na200_1_i;
wire na200_2;
wire na200_2_i;
wire na201_2;
wire na201_2_i;
wire na202_1;
wire na202_1_i;
wire na203_1;
wire na203_2;
wire na204_1;
wire na204_1_i;
wire na204_2;
wire na204_2_i;
wire na205_2;
wire na205_2_i;
wire na207_1;
wire na207_1_i;
wire na207_2;
wire na207_2_i;
wire na208_1;
wire na208_1_i;
wire na209_1;
wire na209_1_i;
wire na210_1;
wire na210_1_i;
wire na211_1;
wire na211_1_i;
wire na212_1;
wire na212_1_i;
wire na214_1;
wire na214_1_i;
wire na214_2;
wire na214_2_i;
wire na216_1;
wire na216_1_i;
wire na216_2;
wire na216_2_i;
wire na217_1;
wire na217_1_i;
wire na217_2;
wire na217_2_i;
wire na218_1;
wire na219_2;
wire na220_1;
wire na221_1;
wire na221_1_i;
wire na222_1;
wire na222_2;
wire na223_2;
wire na224_1;
wire na225_2;
wire na226_1;
wire na226_2;
wire na229_1;
wire na232_1;
wire na232_1_i;
wire na232_2;
wire na232_2_i;
wire na233_1;
wire na233_2;
wire na234_1;
wire na235_2;
wire na236_1;
wire na237_1;
wire na237_1_i;
wire na238_1;
wire na238_1_i;
wire na239_1;
wire na239_1_i;
wire na240_1;
wire na240_1_i;
wire na241_1;
wire na241_1_i;
wire na242_1;
wire na242_1_i;
wire na243_1;
wire na243_1_i;
wire na244_1;
wire na244_1_i;
wire na245_1;
wire na245_1_i;
wire na246_1;
wire na246_1_i;
wire na247_1;
wire na247_1_i;
wire na248_1;
wire na249_1;
wire na251_2;
wire na252_1;
wire na253_1;
wire na254_1;
wire na255_2;
wire na260_2;
wire na261_2;
wire na262_1;
wire na264_1;
wire na264_1_i;
wire na265_1;
wire na265_1_i;
wire na265_2;
wire na265_2_i;
wire na266_1;
wire na266_1_i;
wire na268_1;
wire na268_1_i;
wire na268_2;
wire na268_2_i;
wire na269_2;
wire na269_2_i;
wire na270_1;
wire na270_1_i;
wire na270_2;
wire na270_2_i;
wire na272_1;
wire na272_1_i;
wire na273_1;
wire na273_2;
wire na274_1;
wire na274_1_i;
wire na274_2;
wire na274_2_i;
wire na275_2;
wire na276_1;
wire na277_1;
wire na277_1_i;
wire na280_1;
wire na280_1_i;
wire na280_2;
wire na280_2_i;
wire na281_1;
wire na281_1_i;
wire na281_2;
wire na281_2_i;
wire na282_1;
wire na282_1_i;
wire na283_1;
wire na283_1_i;
wire na284_1;
wire na284_1_i;
wire na285_1;
wire na285_1_i;
wire na285_2;
wire na285_2_i;
wire na287_1;
wire na287_1_i;
wire na287_2;
wire na287_2_i;
wire na288_1;
wire na288_1_i;
wire na288_2;
wire na288_2_i;
wire na289_1;
wire na289_1_i;
wire na292_1;
wire na292_1_i;
wire na292_2;
wire na292_2_i;
wire na293_2;
wire na293_2_i;
wire na294_2;
wire na294_2_i;
wire na295_1;
wire na295_1_i;
wire na295_2;
wire na295_2_i;
wire na297_1;
wire na297_1_i;
wire na297_2;
wire na297_2_i;
wire na299_1;
wire na299_1_i;
wire na301_1;
wire na302_1;
wire na303_2;
wire na304_1;
wire na304_2;
wire na307_1;
wire na310_1;
wire na310_2;
wire na311_1;
wire na311_1_i;
wire na312_1;
wire na312_1_i;
wire na313_1;
wire na313_1_i;
wire na314_1;
wire na314_1_i;
wire na315_1;
wire na315_1_i;
wire na316_1;
wire na316_1_i;
wire na317_2;
wire na318_1;
wire na319_2;
wire na321_1;
wire na322_1;
wire na322_1_i;
wire na323_1;
wire na323_1_i;
wire na324_1;
wire na324_1_i;
wire na325_1;
wire na325_1_i;
wire na326_1;
wire na326_1_i;
wire na327_1;
wire na327_1_i;
wire na328_1;
wire na328_1_i;
wire na329_1;
wire na329_1_i;
wire na330_1;
wire na330_1_i;
wire na331_1;
wire na331_1_i;
wire na332_1;
wire na332_1_i;
wire na333_1;
wire na333_1_i;
wire na335_1;
wire na335_2;
wire na336_2;
wire na337_2;
wire na338_2;
wire na340_2;
wire na341_1;
wire na341_2;
wire na343_1;
wire na346_1;
wire na346_2;
wire na349_2;
wire na349_2_i;
wire na350_1;
wire na351_1;
wire na352_1;
wire na352_2;
wire na353_1;
wire na354_1;
wire na355_1;
wire na356_1;
wire na357_1;
wire na358_2;
wire na358_2_i;
wire na360_1;
wire na360_1_i;
wire na360_2;
wire na360_2_i;
wire na361_1;
wire na361_1_i;
wire na362_1;
wire na362_2;
wire na363_1;
wire na363_2;
wire na364_1;
wire na364_2;
wire na365_1;
wire na365_2;
wire na366_1;
wire na366_2;
wire na367_1;
wire na367_2;
wire na368_1;
wire na368_2;
wire na369_1;
wire na369_2;
wire na370_1;
wire na370_1_i;
wire na371_1;
wire na371_1_i;
wire na372_1;
wire na373_1;
wire na373_1_i;
wire na374_1;
wire na374_1_i;
wire na375_1;
wire na375_1_i;
wire na376_1;
wire na377_1;
wire na377_1_i;
wire na378_1;
wire na378_1_i;
wire na379_1;
wire na379_1_i;
wire na380_1;
wire na380_1_i;
wire na381_1;
wire na381_1_i;
wire na382_1;
wire na382_1_i;
wire na383_1;
wire na383_1_i;
wire na384_1;
wire na384_1_i;
wire na387_2;
wire na387_2_i;
wire na388_1;
wire na388_1_i;
wire na388_2;
wire na388_2_i;
wire na390_1;
wire na390_1_i;
wire na390_2;
wire na390_2_i;
wire na391_1;
wire na391_1_i;
wire na391_2;
wire na391_2_i;
wire na392_1;
wire na392_1_i;
wire na394_1;
wire na395_2;
wire na396_1;
wire na396_1_i;
wire na397_1;
wire na397_1_i;
wire na398_1;
wire na398_1_i;
wire na399_1;
wire na399_2;
wire na402_2;
wire na402_2_i;
wire na403_1;
wire na403_1_i;
wire na403_2;
wire na403_2_i;
wire na405_2;
wire na407_2;
wire na408_1;
wire na409_1;
wire na409_1_i;
wire na410_1;
wire na410_1_i;
wire na411_1;
wire na411_1_i;
wire na412_1;
wire na412_1_i;
wire na413_1;
wire na413_1_i;
wire na414_1;
wire na414_1_i;
wire na415_1;
wire na415_1_i;
wire na416_1;
wire na416_1_i;
wire na417_1;
wire na417_1_i;
wire na418_1;
wire na418_1_i;
wire na420_2;
wire na421_1;
wire na423_1;
wire na423_2;
wire na424_2;
wire na425_2;
wire na426_1;
wire na426_1_i;
wire na427_1;
wire na427_2;
wire na428_1;
wire na428_1_i;
wire na429_1;
wire na429_1_i;
wire na430_2;
wire na430_2_i;
wire na432_2;
wire na432_2_i;
wire na434_1;
wire na434_1_i;
wire na434_2;
wire na434_2_i;
wire na435_1;
wire na435_1_i;
wire na435_2;
wire na435_2_i;
wire na436_1;
wire na437_1;
wire na437_1_i;
wire na438_1;
wire na438_1_i;
wire na439_1;
wire na439_1_i;
wire na440_1;
wire na440_1_i;
wire na441_1;
wire na441_1_i;
wire na442_1;
wire na442_1_i;
wire na443_1;
wire na443_1_i;
wire na445_1;
wire na445_2;
wire na446_2;
wire na447_2;
wire na449_2;
wire na450_1;
wire na450_2;
wire na452_1;
wire na455_1;
wire na455_2;
wire na456_1;
wire na456_1_i;
wire na456_2;
wire na456_2_i;
wire na457_1;
wire na457_1_i;
wire na458_1;
wire na459_1;
wire na460_1;
wire na460_2;
wire na461_1;
wire na462_1;
wire na463_1;
wire na465_1;
wire na466_1;
wire na467_1;
wire na468_2;
wire na469_2;
wire na469_2_i;
wire na470_1;
wire na470_1_i;
wire na471_1;
wire na471_1_i;
wire na472_1;
wire na472_1_i;
wire na473_1;
wire na473_1_i;
wire na474_1;
wire na474_1_i;
wire na475_1;
wire na475_1_i;
wire na476_1;
wire na476_1_i;
wire na477_1;
wire na477_1_i;
wire na478_1;
wire na478_1_i;
wire na479_1;
wire na479_1_i;
wire na480_1;
wire na480_1_i;
wire na481_1;
wire na481_1_i;
wire na482_1;
wire na482_1_i;
wire na483_1;
wire na483_1_i;
wire na484_1;
wire na484_1_i;
wire na485_1;
wire na485_1_i;
wire na486_1;
wire na486_1_i;
wire na487_1;
wire na487_1_i;
wire na488_1;
wire na488_1_i;
wire na489_1;
wire na489_1_i;
wire na490_1;
wire na490_1_i;
wire na491_1;
wire na491_1_i;
wire na492_1;
wire na492_1_i;
wire na493_1;
wire na493_1_i;
wire na494_1;
wire na494_1_i;
wire na495_1;
wire na496_1;
wire na496_1_i;
wire na497_1;
wire na498_1;
wire na499_1;
wire na499_1_i;
wire na500_1;
wire na501_1;
wire na501_1_i;
wire na502_1;
wire na503_1;
wire na503_1_i;
wire na504_1;
wire na505_1;
wire na505_1_i;
wire na506_2;
wire na506_2_i;
wire na507_1;
wire na507_1_i;
wire na508_2;
wire na508_2_i;
wire na510_1;
wire na510_1_i;
wire na511_1;
wire na511_2;
wire na512_1;
wire na513_1;
wire na514_2;
wire na516_1;
wire na517_2;
wire na518_1;
wire na518_1_i;
wire na519_1;
wire na519_2;
wire na520_2;
wire na521_1;
wire na522_2;
wire na523_1;
wire na524_1;
wire na525_1;
wire na525_1_i;
wire na526_1;
wire na528_1;
wire na529_2;
wire na529_2_i;
wire na530_1;
wire na530_2;
wire na531_1;
wire na531_1_i;
wire na532_1;
wire na532_1_i;
wire na533_1;
wire na533_1_i;
wire na534_1;
wire na534_1_i;
wire na534_2;
wire na534_2_i;
wire na535_1;
wire na535_1_i;
wire na536_1;
wire na536_2;
wire na537_1;
wire na537_1_i;
wire na538_1;
wire na538_1_i;
wire na539_1;
wire na539_1_i;
wire na540_1;
wire na540_1_i;
wire na541_1;
wire na541_1_i;
wire na542_1;
wire na542_1_i;
wire na543_1;
wire na543_1_i;
wire na543_2;
wire na543_2_i;
wire na545_1;
wire na545_1_i;
wire na545_2;
wire na545_2_i;
wire na547_1;
wire na547_1_i;
wire na547_2;
wire na547_2_i;
wire na549_1;
wire na549_1_i;
wire na549_2;
wire na549_2_i;
wire na551_1;
wire na551_1_i;
wire na551_2;
wire na551_2_i;
wire na553_1;
wire na553_1_i;
wire na553_2;
wire na553_2_i;
wire na555_1;
wire na555_1_i;
wire na555_2;
wire na555_2_i;
wire na557_1;
wire na557_1_i;
wire na557_2;
wire na557_2_i;
wire na559_1;
wire na559_1_i;
wire na559_2;
wire na559_2_i;
wire na561_1;
wire na561_1_i;
wire na561_2;
wire na561_2_i;
wire na563_1;
wire na563_1_i;
wire na563_2;
wire na563_2_i;
wire na565_1;
wire na565_1_i;
wire na565_2;
wire na565_2_i;
wire na567_1;
wire na567_1_i;
wire na567_2;
wire na567_2_i;
wire na569_1;
wire na569_1_i;
wire na569_2;
wire na569_2_i;
wire na571_1;
wire na571_1_i;
wire na571_2;
wire na571_2_i;
wire na573_1;
wire na573_1_i;
wire na573_2;
wire na573_2_i;
wire na575_1;
wire na576_2;
wire na576_2_i;
wire na577_1;
wire na578_1;
wire na578_1_i;
wire na579_1;
wire na579_1_i;
wire na580_1;
wire na580_1_i;
wire na582_2;
wire na582_2_i;
wire na584_1;
wire na584_1_i;
wire na586_1;
wire na586_1_i;
wire na588_1;
wire na588_1_i;
wire na590_1;
wire na590_1_i;
wire na591_1;
wire na591_1_i;
wire na592_1;
wire na592_1_i;
wire na593_1;
wire na593_1_i;
wire na594_1;
wire na594_1_i;
wire na595_1;
wire na595_1_i;
wire na596_1;
wire na596_1_i;
wire na597_1;
wire na597_2;
wire na598_1;
wire na598_2;
wire na599_2;
wire na600_2;
wire na603_1;
wire na603_2;
wire na605_1;
wire na606_1;
wire na607_1;
wire na612_1;
wire na613_2;
wire na614_1;
wire na618_1;
wire na619_1;
wire na620_1;
wire na620_1_i;
wire na621_1;
wire na622_1;
wire na623_2;
wire na624_1;
wire na625_2;
wire na626_1;
wire na627_1;
wire na628_1;
wire na629_1;
wire na630_1;
wire na631_2;
wire na632_1;
wire na633_1;
wire na633_1_i;
wire na634_1;
wire na634_1_i;
wire na635_1;
wire na635_1_i;
wire na636_1;
wire na638_2;
wire na638_2_i;
wire na639_1;
wire na639_2;
wire na640_1;
wire na640_1_i;
wire na641_1;
wire na641_1_i;
wire na642_1;
wire na642_1_i;
wire na643_2;
wire na644_1;
wire na645_1;
wire na645_1_i;
wire na647_1;
wire na647_1_i;
wire na648_1;
wire na648_1_i;
wire na649_1;
wire na649_1_i;
wire na650_1;
wire na650_1_i;
wire na651_1;
wire na651_1_i;
wire na652_1;
wire na652_1_i;
wire na653_1;
wire na653_1_i;
wire na654_1;
wire na654_1_i;
wire na655_1;
wire na655_1_i;
wire na656_1;
wire na656_1_i;
wire na657_1;
wire na657_1_i;
wire na658_1;
wire na658_1_i;
wire na659_1;
wire na659_1_i;
wire na660_1;
wire na660_1_i;
wire na661_1;
wire na661_1_i;
wire na662_1;
wire na662_1_i;
wire na663_1;
wire na663_1_i;
wire na664_1;
wire na664_1_i;
wire na665_1;
wire na665_1_i;
wire na666_1;
wire na666_1_i;
wire na667_1;
wire na667_1_i;
wire na668_1;
wire na668_1_i;
wire na669_1;
wire na669_1_i;
wire na670_1;
wire na670_1_i;
wire na671_1;
wire na671_1_i;
wire na672_1;
wire na672_1_i;
wire na673_1;
wire na674_1;
wire na674_1_i;
wire na675_1;
wire na675_1_i;
wire na676_1;
wire na677_2;
wire na678_1;
wire na678_1_i;
wire na679_1;
wire na680_1;
wire na680_1_i;
wire na681_1;
wire na682_1;
wire na682_1_i;
wire na683_1;
wire na684_1;
wire na684_1_i;
wire na685_1;
wire na685_1_i;
wire na686_1;
wire na686_1_i;
wire na687_2;
wire na688_1;
wire na689_1;
wire na690_1;
wire na690_1_i;
wire na692_1;
wire na692_1_i;
wire na693_1;
wire na693_1_i;
wire na694_1;
wire na694_1_i;
wire na695_1;
wire na695_1_i;
wire na696_1;
wire na696_1_i;
wire na697_1;
wire na697_1_i;
wire na698_1;
wire na698_1_i;
wire na699_1;
wire na699_1_i;
wire na700_1;
wire na700_1_i;
wire na701_1;
wire na701_1_i;
wire na702_1;
wire na702_1_i;
wire na703_1;
wire na703_1_i;
wire na704_1;
wire na704_2;
wire na705_1;
wire na706_1;
wire na707_1;
wire na708_2;
wire na709_1;
wire na709_1_i;
wire na710_1;
wire na710_1_i;
wire na711_1;
wire na711_1_i;
wire na712_1;
wire na712_1_i;
wire na713_1;
wire na713_1_i;
wire na713_2;
wire na713_2_i;
wire na714_1;
wire na714_1_i;
wire na715_1;
wire na715_1_i;
wire na716_1;
wire na716_1_i;
wire na717_1;
wire na717_1_i;
wire na718_1;
wire na718_1_i;
wire na719_1;
wire na719_1_i;
wire na720_1;
wire na720_1_i;
wire na721_1;
wire na721_1_i;
wire na722_1;
wire na722_1_i;
wire na723_1;
wire na723_1_i;
wire na724_1;
wire na724_1_i;
wire na725_1;
wire na725_1_i;
wire na726_1;
wire na726_1_i;
wire na727_1;
wire na727_1_i;
wire na728_1;
wire na728_1_i;
wire na728_2;
wire na728_2_i;
wire na730_1;
wire na730_1_i;
wire na730_2;
wire na730_2_i;
wire na732_1;
wire na732_1_i;
wire na732_2;
wire na732_2_i;
wire na734_1;
wire na734_1_i;
wire na734_2;
wire na734_2_i;
wire na736_1;
wire na736_1_i;
wire na736_2;
wire na736_2_i;
wire na738_1;
wire na738_1_i;
wire na738_2;
wire na738_2_i;
wire na740_1;
wire na740_1_i;
wire na740_2;
wire na740_2_i;
wire na742_1;
wire na742_1_i;
wire na742_2;
wire na742_2_i;
wire na744_1;
wire na744_1_i;
wire na744_2;
wire na744_2_i;
wire na746_1;
wire na746_1_i;
wire na746_2;
wire na746_2_i;
wire na748_1;
wire na748_1_i;
wire na748_2;
wire na748_2_i;
wire na750_1;
wire na750_1_i;
wire na750_2;
wire na750_2_i;
wire na752_1;
wire na752_1_i;
wire na752_2;
wire na752_2_i;
wire na754_1;
wire na754_1_i;
wire na754_2;
wire na754_2_i;
wire na756_1;
wire na756_1_i;
wire na756_2;
wire na756_2_i;
wire na758_1;
wire na758_1_i;
wire na758_2;
wire na758_2_i;
wire na760_1;
wire na760_1_i;
wire na761_2;
wire na762_1;
wire na762_1_i;
wire na763_2;
wire na763_2_i;
wire na764_1;
wire na765_1;
wire na765_1_i;
wire na766_1;
wire na766_1_i;
wire na767_1;
wire na767_1_i;
wire na769_1;
wire na769_1_i;
wire na771_2;
wire na771_2_i;
wire na773_2;
wire na773_2_i;
wire na775_2;
wire na775_2_i;
wire na777_1;
wire na777_1_i;
wire na778_1;
wire na778_1_i;
wire na779_1;
wire na779_1_i;
wire na780_1;
wire na780_1_i;
wire na781_1;
wire na781_1_i;
wire na782_1;
wire na782_1_i;
wire na783_1;
wire na783_1_i;
wire na784_1;
wire na784_2;
wire na785_1;
wire na785_2;
wire na786_1;
wire na787_1;
wire na790_1;
wire na790_2;
wire na792_1;
wire na796_2;
wire na797_1;
wire na798_1;
wire na798_1_i;
wire na799_1;
wire na800_1;
wire na801_2;
wire na802_1;
wire na803_1;
wire na804_1;
wire na805_1;
wire na806_1;
wire na807_2;
wire na808_1;
wire na809_1;
wire na810_1;
wire na811_1;
wire na811_1_i;
wire na812_1;
wire na813_1;
wire na814_1;
wire na814_1_i;
wire na815_1;
wire na815_1_i;
wire na816_1;
wire na816_1_i;
wire na817_1;
wire na819_2;
wire na820_1;
wire na821_1;
wire na821_1_i;
wire na822_1;
wire na822_2;
wire na823_1;
wire na823_1_i;
wire na825_1;
wire na825_1_i;
wire na826_1;
wire na826_1_i;
wire na826_2;
wire na826_2_i;
wire na827_1;
wire na827_1_i;
wire na828_1;
wire na828_1_i;
wire na829_1;
wire na829_1_i;
wire na830_1;
wire na830_1_i;
wire na831_1;
wire na831_1_i;
wire na832_1;
wire na832_1_i;
wire na833_1;
wire na833_1_i;
wire na834_1;
wire na834_1_i;
wire na835_1;
wire na835_1_i;
wire na836_1;
wire na836_1_i;
wire na837_1;
wire na837_1_i;
wire na838_1;
wire na838_1_i;
wire na839_1;
wire na839_1_i;
wire na840_1;
wire na840_1_i;
wire na841_1;
wire na841_1_i;
wire na842_1;
wire na842_1_i;
wire na843_1;
wire na843_1_i;
wire na844_1;
wire na844_1_i;
wire na845_1;
wire na845_1_i;
wire na846_1;
wire na846_1_i;
wire na847_1;
wire na847_1_i;
wire na848_1;
wire na848_1_i;
wire na849_1;
wire na849_1_i;
wire na850_1;
wire na850_1_i;
wire na851_1;
wire na851_1_i;
wire na852_1;
wire na853_1;
wire na853_1_i;
wire na854_1;
wire na855_1;
wire na856_1;
wire na856_1_i;
wire na857_1;
wire na858_1;
wire na858_1_i;
wire na859_1;
wire na860_1;
wire na860_1_i;
wire na861_1;
wire na862_1;
wire na862_1_i;
wire na864_1;
wire na864_1_i;
wire na865_1;
wire na865_1_i;
wire na866_1;
wire na866_1_i;
wire na867_1;
wire na867_1_i;
wire na868_1;
wire na868_1_i;
wire na869_1;
wire na869_1_i;
wire na870_1;
wire na870_1_i;
wire na871_1;
wire na871_1_i;
wire na872_1;
wire na872_1_i;
wire na873_1;
wire na873_1_i;
wire na874_1;
wire na874_1_i;
wire na875_1;
wire na875_1_i;
wire na876_1;
wire na876_1_i;
wire na877_1;
wire na877_2;
wire na878_1;
wire na879_1;
wire na880_2;
wire na881_1;
wire na881_2;
wire na882_2;
wire na883_1;
wire na884_2;
wire na885_1;
wire na886_1;
wire na886_1_i;
wire na887_2;
wire na887_2_i;
wire na888_1;
wire na888_2;
wire na891_1;
wire na891_1_i;
wire na891_2;
wire na891_2_i;
wire na892_1;
wire na892_1_i;
wire na892_2;
wire na892_2_i;
wire na894_1;
wire na894_1_i;
wire na894_2;
wire na894_2_i;
wire na896_1;
wire na896_1_i;
wire na896_2;
wire na896_2_i;
wire na898_1;
wire na898_1_i;
wire na898_2;
wire na898_2_i;
wire na900_1;
wire na900_1_i;
wire na900_2;
wire na900_2_i;
wire na902_1;
wire na902_1_i;
wire na902_2;
wire na902_2_i;
wire na904_1;
wire na904_1_i;
wire na904_2;
wire na904_2_i;
wire na906_1;
wire na906_1_i;
wire na906_2;
wire na906_2_i;
wire na908_1;
wire na908_1_i;
wire na908_2;
wire na908_2_i;
wire na910_1;
wire na910_1_i;
wire na910_2;
wire na910_2_i;
wire na912_1;
wire na912_1_i;
wire na912_2;
wire na912_2_i;
wire na914_1;
wire na914_1_i;
wire na914_2;
wire na914_2_i;
wire na916_1;
wire na916_1_i;
wire na916_2;
wire na916_2_i;
wire na918_1;
wire na918_1_i;
wire na918_2;
wire na918_2_i;
wire na920_1;
wire na920_1_i;
wire na920_2;
wire na920_2_i;
wire na922_1;
wire na922_1_i;
wire na922_2;
wire na922_2_i;
wire na924_1;
wire na926_1;
wire na926_1_i;
wire na927_1;
wire na927_1_i;
wire na927_2;
wire na927_2_i;
wire na928_1;
wire na928_1_i;
wire na929_1;
wire na929_1_i;
wire na930_2;
wire na930_2_i;
wire na931_1;
wire na932_1;
wire na932_1_i;
wire na933_1;
wire na933_1_i;
wire na934_1;
wire na934_1_i;
wire na936_2;
wire na936_2_i;
wire na938_1;
wire na938_1_i;
wire na940_2;
wire na940_2_i;
wire na942_1;
wire na942_1_i;
wire na944_1;
wire na944_1_i;
wire na945_1;
wire na945_1_i;
wire na946_1;
wire na946_1_i;
wire na947_1;
wire na947_1_i;
wire na948_1;
wire na948_1_i;
wire na949_1;
wire na949_1_i;
wire na950_1;
wire na950_1_i;
wire na951_1;
wire na951_2;
wire na952_1;
wire na952_2;
wire na953_2;
wire na954_1;
wire na957_1;
wire na957_2;
wire na959_1;
wire na963_2;
wire na964_1;
wire na965_1;
wire na965_1_i;
wire na966_1;
wire na967_1;
wire na968_2;
wire na969_1;
wire na970_2;
wire na971_1;
wire na972_2;
wire na973_1;
wire na974_1;
wire na975_1;
wire na976_2;
wire na977_1;
wire na978_1;
wire na978_1_i;
wire na980_2;
wire na980_2_i;
wire na982_2;
wire na983_2;
wire na984_1;
wire na984_1_i;
wire na986_1;
wire na986_1_i;
wire na986_2;
wire na986_2_i;
wire na987_1;
wire na987_1_i;
wire na990_1;
wire na992_1;
wire na993_1;
wire na993_1_i;
wire na994_1;
wire na994_1_i;
wire na995_1;
wire na995_1_i;
wire na996_1;
wire na996_1_i;
wire na997_1;
wire na997_1_i;
wire na998_1;
wire na998_1_i;
wire na999_1;
wire na999_1_i;
wire na1000_1;
wire na1000_1_i;
wire na1001_1;
wire na1001_1_i;
wire na1002_1;
wire na1002_1_i;
wire na1003_1;
wire na1003_1_i;
wire na1004_1;
wire na1004_1_i;
wire na1005_1;
wire na1005_1_i;
wire na1006_1;
wire na1006_1_i;
wire na1007_1;
wire na1007_1_i;
wire na1008_1;
wire na1008_1_i;
wire na1009_1;
wire na1009_1_i;
wire na1010_1;
wire na1010_1_i;
wire na1011_1;
wire na1011_1_i;
wire na1012_1;
wire na1012_1_i;
wire na1013_1;
wire na1013_1_i;
wire na1014_1;
wire na1014_1_i;
wire na1015_1;
wire na1015_1_i;
wire na1016_1;
wire na1016_1_i;
wire na1017_1;
wire na1017_1_i;
wire na1018_1;
wire na1018_1_i;
wire na1019_1;
wire na1019_1_i;
wire na1020_1;
wire na1020_1_i;
wire na1021_1;
wire na1021_1_i;
wire na1022_1;
wire na1022_1_i;
wire na1023_1;
wire na1023_1_i;
wire na1024_1;
wire na1024_1_i;
wire na1025_1;
wire na1026_1;
wire na1026_1_i;
wire na1027_1;
wire na1028_1;
wire na1029_1;
wire na1029_1_i;
wire na1030_1;
wire na1031_1;
wire na1031_1_i;
wire na1032_1;
wire na1033_1;
wire na1033_1_i;
wire na1034_1;
wire na1035_1;
wire na1035_1_i;
wire na1036_1;
wire na1036_1_i;
wire na1037_1;
wire na1037_2;
wire na1038_1;
wire na1039_1;
wire na1040_2;
wire na1042_1;
wire na1043_1;
wire na1044_1;
wire na1044_2;
wire na1045_2;
wire na1046_1;
wire na1047_1;
wire na1048_1;
wire na1049_1;
wire na1050_1;
wire na1050_1_i;
wire na1051_1;
wire na1051_1_i;
wire na1051_2;
wire na1051_2_i;
wire na1052_1;
wire na1052_1_i;
wire na1052_2;
wire na1052_2_i;
wire na1054_1;
wire na1054_1_i;
wire na1054_2;
wire na1054_2_i;
wire na1056_1;
wire na1056_1_i;
wire na1056_2;
wire na1056_2_i;
wire na1058_1;
wire na1058_1_i;
wire na1058_2;
wire na1058_2_i;
wire na1060_1;
wire na1060_1_i;
wire na1060_2;
wire na1060_2_i;
wire na1062_1;
wire na1062_1_i;
wire na1062_2;
wire na1062_2_i;
wire na1064_1;
wire na1064_1_i;
wire na1064_2;
wire na1064_2_i;
wire na1066_1;
wire na1066_1_i;
wire na1066_2;
wire na1066_2_i;
wire na1068_1;
wire na1068_1_i;
wire na1068_2;
wire na1068_2_i;
wire na1070_1;
wire na1070_1_i;
wire na1070_2;
wire na1070_2_i;
wire na1072_1;
wire na1072_1_i;
wire na1072_2;
wire na1072_2_i;
wire na1074_1;
wire na1074_1_i;
wire na1074_2;
wire na1074_2_i;
wire na1076_1;
wire na1076_1_i;
wire na1076_2;
wire na1076_2_i;
wire na1078_1;
wire na1078_1_i;
wire na1078_2;
wire na1078_2_i;
wire na1080_1;
wire na1080_1_i;
wire na1080_2;
wire na1080_2_i;
wire na1082_1;
wire na1082_1_i;
wire na1082_2;
wire na1082_2_i;
wire na1084_2;
wire na1085_1;
wire na1085_1_i;
wire na1086_1;
wire na1087_1;
wire na1088_1;
wire na1089_2;
wire na1090_1;
wire na1090_1_i;
wire na1091_2;
wire na1091_2_i;
wire na1092_1;
wire na1093_1;
wire na1093_1_i;
wire na1094_1;
wire na1094_1_i;
wire na1095_1;
wire na1095_1_i;
wire na1097_2;
wire na1097_2_i;
wire na1099_2;
wire na1099_2_i;
wire na1101_2;
wire na1101_2_i;
wire na1103_1;
wire na1103_1_i;
wire na1105_1;
wire na1105_1_i;
wire na1106_1;
wire na1106_1_i;
wire na1107_1;
wire na1107_1_i;
wire na1108_1;
wire na1108_1_i;
wire na1109_1;
wire na1109_1_i;
wire na1110_1;
wire na1110_1_i;
wire na1111_1;
wire na1111_1_i;
wire na1112_1;
wire na1112_2;
wire na1113_1;
wire na1113_2;
wire na1114_1;
wire na1115_2;
wire na1118_1;
wire na1118_2;
wire na1120_2;
wire na1121_1;
wire na1122_2;
wire na1127_2;
wire na1128_2;
wire na1129_1;
wire na1133_1;
wire na1134_1;
wire na1135_1;
wire na1135_1_i;
wire na1136_1;
wire na1137_1;
wire na1138_1;
wire na1139_1;
wire na1140_1;
wire na1141_1;
wire na1142_2;
wire na1143_1;
wire na1144_2;
wire na1145_1;
wire na1146_1;
wire na1147_1;
wire na1148_2;
wire na1149_1;
wire na1149_1_i;
wire na1149_2;
wire na1149_2_i;
wire na1151_1;
wire na1151_1_i;
wire na1152_1;
wire na1152_1_i;
wire na1153_1;
wire na1153_1_i;
wire na1154_1;
wire na1154_1_i;
wire na1155_1;
wire na1155_1_i;
wire na1156_1;
wire na1156_1_i;
wire na1157_1;
wire na1157_1_i;
wire na1158_1;
wire na1158_1_i;
wire na1159_1;
wire na1159_1_i;
wire na1160_1;
wire na1160_1_i;
wire na1161_1;
wire na1161_1_i;
wire na1162_1;
wire na1162_1_i;
wire na1163_1;
wire na1163_1_i;
wire na1164_1;
wire na1164_1_i;
wire na1165_1;
wire na1165_1_i;
wire na1166_1;
wire na1166_1_i;
wire na1167_1;
wire na1167_1_i;
wire na1168_1;
wire na1168_1_i;
wire na1169_1;
wire na1169_1_i;
wire na1170_1;
wire na1170_1_i;
wire na1171_1;
wire na1171_1_i;
wire na1172_1;
wire na1172_1_i;
wire na1173_1;
wire na1173_1_i;
wire na1174_1;
wire na1174_1_i;
wire na1175_1;
wire na1175_1_i;
wire na1176_1;
wire na1177_1;
wire na1177_1_i;
wire na1178_1;
wire na1179_1;
wire na1180_1;
wire na1180_1_i;
wire na1181_1;
wire na1182_1;
wire na1182_1_i;
wire na1183_1;
wire na1184_1;
wire na1184_1_i;
wire na1185_1;
wire na1186_1;
wire na1186_1_i;
wire na1187_1;
wire na1187_1_i;
wire na1188_1;
wire na1188_1_i;
wire na1191_1;
wire na1192_1;
wire na1192_2;
wire na1193_1;
wire na1194_1;
wire na1195_2;
wire na1196_1;
wire na1197_1;
wire na1198_1;
wire na1198_1_i;
wire na1199_1;
wire na1199_1_i;
wire na1199_2;
wire na1199_2_i;
wire na1200_1;
wire na1200_1_i;
wire na1200_2;
wire na1200_2_i;
wire na1202_1;
wire na1202_1_i;
wire na1202_2;
wire na1202_2_i;
wire na1204_1;
wire na1204_1_i;
wire na1204_2;
wire na1204_2_i;
wire na1206_1;
wire na1206_1_i;
wire na1206_2;
wire na1206_2_i;
wire na1208_1;
wire na1208_1_i;
wire na1208_2;
wire na1208_2_i;
wire na1210_1;
wire na1210_1_i;
wire na1210_2;
wire na1210_2_i;
wire na1212_1;
wire na1212_1_i;
wire na1212_2;
wire na1212_2_i;
wire na1214_1;
wire na1214_1_i;
wire na1214_2;
wire na1214_2_i;
wire na1216_1;
wire na1216_1_i;
wire na1216_2;
wire na1216_2_i;
wire na1218_1;
wire na1218_1_i;
wire na1218_2;
wire na1218_2_i;
wire na1220_1;
wire na1220_1_i;
wire na1220_2;
wire na1220_2_i;
wire na1222_1;
wire na1222_1_i;
wire na1222_2;
wire na1222_2_i;
wire na1224_1;
wire na1224_1_i;
wire na1224_2;
wire na1224_2_i;
wire na1226_1;
wire na1226_1_i;
wire na1226_2;
wire na1226_2_i;
wire na1228_1;
wire na1228_1_i;
wire na1228_2;
wire na1228_2_i;
wire na1230_1;
wire na1230_1_i;
wire na1230_2;
wire na1230_2_i;
wire na1232_2;
wire na1233_1;
wire na1233_1_i;
wire na1234_1;
wire na1235_1;
wire na1235_1_i;
wire na1236_1;
wire na1236_1_i;
wire na1237_2;
wire na1237_2_i;
wire na1239_1;
wire na1239_1_i;
wire na1241_2;
wire na1241_2_i;
wire na1243_1;
wire na1243_1_i;
wire na1245_1;
wire na1245_1_i;
wire na1247_1;
wire na1247_1_i;
wire na1248_1;
wire na1248_1_i;
wire na1249_1;
wire na1249_1_i;
wire na1250_1;
wire na1250_1_i;
wire na1251_1;
wire na1251_1_i;
wire na1252_1;
wire na1252_1_i;
wire na1253_1;
wire na1253_1_i;
wire na1254_1;
wire na1254_2;
wire na1255_1;
wire na1255_2;
wire na1256_2;
wire na1257_1;
wire na1260_1;
wire na1260_2;
wire na1262_1;
wire na1263_1;
wire na1264_1;
wire na1269_1;
wire na1270_2;
wire na1271_1;
wire na1275_1;
wire na1276_1;
wire na1277_1;
wire na1277_1_i;
wire na1278_1;
wire na1279_1;
wire na1280_1;
wire na1281_1;
wire na1282_2;
wire na1283_1;
wire na1284_2;
wire na1285_1;
wire na1286_2;
wire na1287_1;
wire na1288_1;
wire na1289_1;
wire na1290_1;
wire na1290_1_i;
wire na1292_1;
wire na1292_1_i;
wire na1293_1;
wire na1293_1_i;
wire na1294_1;
wire na1294_1_i;
wire na1295_1;
wire na1295_1_i;
wire na1296_1;
wire na1296_1_i;
wire na1296_2;
wire na1296_2_i;
wire na1297_1;
wire na1298_1;
wire na1298_1_i;
wire na1301_1;
wire na1301_1_i;
wire na1302_1;
wire na1302_1_i;
wire na1303_1;
wire na1303_1_i;
wire na1304_1;
wire na1304_1_i;
wire na1304_2;
wire na1304_2_i;
wire na1305_2;
wire na1305_2_i;
wire na1306_1;
wire na1306_1_i;
wire na1306_2;
wire na1306_2_i;
wire na1307_1;
wire na1307_1_i;
wire na1307_2;
wire na1307_2_i;
wire na1308_1;
wire na1308_1_i;
wire na1309_1;
wire na1309_1_i;
wire na1310_1;
wire na1311_2;
wire na1312_1;
wire na1312_1_i;
wire na1313_1;
wire na1313_1_i;
wire na1314_2;
wire na1314_2_i;
wire na1315_2;
wire na1316_1;
wire na1317_1;
wire na1317_1_i;
wire na1318_1;
wire na1318_1_i;
wire na1319_1;
wire na1319_1_i;
wire na1320_1;
wire na1320_1_i;
wire na1321_1;
wire na1321_1_i;
wire na1322_1;
wire na1322_1_i;
wire na1323_1;
wire na1323_1_i;
wire na1324_1;
wire na1324_1_i;
wire na1325_1;
wire na1325_1_i;
wire na1326_1;
wire na1326_1_i;
wire na1327_1;
wire na1327_1_i;
wire na1328_1;
wire na1328_1_i;
wire na1329_1;
wire na1329_1_i;
wire na1330_1;
wire na1330_1_i;
wire na1330_2;
wire na1330_2_i;
wire na1331_1;
wire na1331_1_i;
wire na1332_1;
wire na1332_1_i;
wire na1333_1;
wire na1334_2;
wire na1335_1;
wire na1335_1_i;
wire na1336_1;
wire na1336_1_i;
wire na1337_1;
wire na1337_1_i;
wire na1338_1;
wire na1338_1_i;
wire na1339_1;
wire na1339_1_i;
wire na1340_1;
wire na1340_1_i;
wire na1341_2;
wire na1341_2_i;
wire na1342_1;
wire na1343_1;
wire na1344_2;
wire na1345_1;
wire na1346_1;
wire na1346_1_i;
wire na1347_1;
wire na1347_1_i;
wire na1349_1;
wire na1349_2;
wire na1350_2;
wire na1350_2_i;
wire na1351_2;
wire na1351_2_i;
wire na1352_1;
wire na1352_1_i;
wire na1353_1;
wire na1353_1_i;
wire na1354_1;
wire na1354_1_i;
wire na1355_1;
wire na1355_1_i;
wire na1356_1;
wire na1356_1_i;
wire na1357_1;
wire na1357_1_i;
wire na1358_1;
wire na1358_1_i;
wire na1359_1;
wire na1359_1_i;
wire na1360_1;
wire na1360_1_i;
wire na1361_1;
wire na1361_1_i;
wire na1362_1;
wire na1362_1_i;
wire na1363_1;
wire na1363_1_i;
wire na1364_1;
wire na1364_1_i;
wire na1365_1;
wire na1365_1_i;
wire na1366_1;
wire na1366_1_i;
wire na1367_1;
wire na1367_1_i;
wire na1368_1;
wire na1368_1_i;
wire na1369_1;
wire na1369_1_i;
wire na1370_2;
wire na1370_2_i;
wire na1371_1;
wire na1372_1;
wire na1373_2;
wire na1374_2;
wire na1375_2;
wire na1375_2_i;
wire na1376_1;
wire na1376_1_i;
wire na1377_1;
wire na1377_1_i;
wire na1378_1;
wire na1378_1_i;
wire na1379_1;
wire na1379_1_i;
wire na1381_1;
wire na1381_1_i;
wire na1383_2;
wire na1383_2_i;
wire na1385_1;
wire na1385_1_i;
wire na1385_2;
wire na1385_2_i;
wire na1386_1;
wire na1386_1_i;
wire na1387_1;
wire na1387_1_i;
wire na1388_1;
wire na1388_1_i;
wire na1389_1;
wire na1389_1_i;
wire na1390_1;
wire na1390_1_i;
wire na1391_1;
wire na1391_1_i;
wire na1392_1;
wire na1392_1_i;
wire na1393_1;
wire na1393_1_i;
wire na1394_1;
wire na1394_1_i;
wire na1395_1;
wire na1395_1_i;
wire na1396_1;
wire na1396_1_i;
wire na1397_1;
wire na1397_1_i;
wire na1398_1;
wire na1399_1;
wire na1400_1;
wire na1401_2;
wire na1402_2;
wire na1403_1;
wire na1404_1;
wire na1405_2;
wire na1406_2;
wire na1407_1;
wire na1408_1;
wire na1409_1;
wire na1410_1;
wire na1411_1;
wire na1412_1;
wire na1413_1;
wire na1414_2;
wire na1415_2;
wire na1416_1;
wire na1417_2;
wire na1418_2;
wire na1419_2;
wire na1420_1;
wire na1421_1;
wire na1422_1;
wire na1423_2;
wire na1424_2;
wire na1425_2;
wire na1426_2;
wire na1427_2;
wire na1428_1;
wire na1429_2;
wire na1431_1;
wire na1432_1;
wire na1432_1_i;
wire na1434_1;
wire na1435_1;
wire na1436_2;
wire na1437_1;
wire na1438_1;
wire na1438_1_i;
wire na1439_1;
wire na1439_1_i;
wire na1440_2;
wire na1440_2_i;
wire na1441_2;
wire na1441_2_i;
wire na1443_1;
wire na1443_1_i;
wire na1443_2;
wire na1443_2_i;
wire na1444_1;
wire na1444_1_i;
wire na1445_1;
wire na1445_2;
wire na1446_2;
wire na1446_2_i;
wire na1447_1;
wire na1447_1_i;
wire na1448_1;
wire na1449_2;
wire na1450_2;
wire na1451_1;
wire na1451_1_i;
wire na1453_2;
wire na1454_2;
wire na1454_2_i;
wire na1456_1;
wire na1457_1;
wire na1458_2;
wire na1459_2;
wire na1460_2;
wire na1460_2_i;
wire na1461_1;
wire na1461_1_i;
wire na1462_2;
wire na1462_2_i;
wire na1463_1;
wire na1463_1_i;
wire na1465_1;
wire na1465_1_i;
wire na1465_2;
wire na1465_2_i;
wire na1466_1;
wire na1466_1_i;
wire na1467_1;
wire na1467_2;
wire na1468_1;
wire na1468_1_i;
wire na1469_1;
wire na1469_1_i;
wire na1470_1;
wire na1471_2;
wire na1472_1;
wire na1473_2;
wire na1473_2_i;
wire na1475_1;
wire na1476_2;
wire na1476_2_i;
wire na1478_1;
wire na1479_1;
wire na1480_1;
wire na1481_2;
wire na1482_2;
wire na1482_2_i;
wire na1483_2;
wire na1483_2_i;
wire na1484_2;
wire na1484_2_i;
wire na1485_1;
wire na1485_1_i;
wire na1487_1;
wire na1487_1_i;
wire na1487_2;
wire na1487_2_i;
wire na1488_1;
wire na1488_1_i;
wire na1489_1;
wire na1489_2;
wire na1490_2;
wire na1490_2_i;
wire na1491_1;
wire na1491_1_i;
wire na1492_1;
wire na1493_2;
wire na1494_2;
wire na1495_2;
wire na1495_2_i;
wire na1497_2;
wire na1498_1;
wire na1498_1_i;
wire na1500_1;
wire na1501_1;
wire na1502_1;
wire na1503_2;
wire na1504_2;
wire na1504_2_i;
wire na1505_2;
wire na1505_2_i;
wire na1506_1;
wire na1506_1_i;
wire na1507_1;
wire na1507_1_i;
wire na1509_2;
wire na1509_2_i;
wire na1510_1;
wire na1510_1_i;
wire na1511_1;
wire na1511_2;
wire na1512_1;
wire na1512_1_i;
wire na1513_1;
wire na1513_1_i;
wire na1514_2;
wire na1515_2;
wire na1516_2;
wire na1517_2;
wire na1517_2_i;
wire na1519_1;
wire na1520_2;
wire na1520_2_i;
wire na1522_1;
wire na1523_1;
wire na1524_2;
wire na1525_1;
wire na1526_1;
wire na1526_1_i;
wire na1527_2;
wire na1527_2_i;
wire na1528_2;
wire na1528_2_i;
wire na1529_2;
wire na1529_2_i;
wire na1531_2;
wire na1531_2_i;
wire na1532_1;
wire na1532_1_i;
wire na1533_1;
wire na1533_2;
wire na1534_2;
wire na1534_2_i;
wire na1535_1;
wire na1535_1_i;
wire na1536_1;
wire na1537_2;
wire na1538_2;
wire na1539_1;
wire na1539_1_i;
wire na1540_2;
wire na1541_1;
wire na1541_1_i;
wire na1541_2;
wire na1541_2_i;
wire na1542_1;
wire na1542_1_i;
wire na1542_2;
wire na1542_2_i;
wire na1543_1;
wire na1543_1_i;
wire na1543_2;
wire na1543_2_i;
wire na1544_1;
wire na1544_1_i;
wire na1544_2;
wire na1544_2_i;
wire na1545_1;
wire na1545_1_i;
wire na1545_2;
wire na1545_2_i;
wire na1564_1;
wire na1567_1;
wire na1567_2;
wire na1570_1;
wire na1574_1;
wire na1576_1;
wire na1577_1;
wire na1578_1;
wire na1579_1;
wire na1579_1_i;
wire na1580_1;
wire na1581_1;
wire na1581_2;
wire na1582_1;
wire na1583_1;
wire na1584_1;
wire na1585_1;
wire na1585_1_i;
wire na1586_1;
wire na1587_1;
wire na1587_2;
wire na1588_1;
wire na1589_1;
wire na1590_1;
wire na1591_1;
wire na1591_1_i;
wire na1592_1;
wire na1593_1;
wire na1593_2;
wire na1594_1;
wire na1595_1;
wire na1596_1;
wire na1597_1;
wire na1597_1_i;
wire na1598_1;
wire na1599_1;
wire na1599_2;
wire na1600_1;
wire na1601_1;
wire na1602_1;
wire na1603_1;
wire na1603_1_i;
wire na1604_1;
wire na1605_1;
wire na1605_2;
wire na1608_1;
wire na1610_1;
wire na1610_2;
wire na1610_4;
wire na1612_1;
wire na1612_4;
wire na1613_1;
wire na1614_1;
wire na1614_2;
wire na1614_4;
wire na1616_1;
wire na1616_4;
wire na1617_1;
wire na1618_1;
wire na1618_2;
wire na1618_4;
wire na1620_1;
wire na1620_2;
wire na1620_4;
wire na1622_1;
wire na1622_2;
wire na1622_4;
wire na1624_1;
wire na1624_2;
wire na1624_4;
wire na1626_1;
wire na1627_1;
wire na1627_4;
wire na1628_1;
wire na1628_2;
wire na1628_4;
wire na1630_1;
wire na1630_2;
wire na1632_1;
wire na1632_4;
wire na1633_1;
wire na1633_2;
wire na1633_4;
wire na1635_1;
wire na1635_2;
wire na1635_4;
wire na1637_1;
wire na1638_1;
wire na1638_4;
wire na1639_1;
wire na1639_2;
wire na1639_4;
wire na1641_1;
wire na1641_2;
wire na1643_1;
wire na1643_2;
wire na1643_4;
wire na1645_1;
wire na1646_4;
wire na1648_1;
wire na1648_4;
wire na1649_1;
wire na1649_2;
wire na1649_4;
wire na1651_1;
wire na1652_1;
wire na1652_4;
wire na1653_1;
wire na1653_2;
wire na1653_4;
wire na1655_1;
wire na1655_2;
wire na1657_1;
wire na1657_4;
wire na1658_1;
wire na1658_2;
wire na1658_4;
wire na1660_1;
wire na1660_2;
wire na1662_4;
wire na1664_1;
wire na1664_4;
wire na1665_1;
wire na1665_4;
wire na1666_1;
wire na1666_2;
wire na1666_4;
wire na1668_1;
wire na1668_2;
wire na1668_4;
wire na1670_1;
wire na1671_4;
wire na1673_1;
wire na1673_4;
wire na1674_1;
wire na1674_2;
wire na1674_4;
wire na1676_1;
wire na1677_1;
wire na1677_4;
wire na1678_1;
wire na1678_2;
wire na1678_4;
wire na1680_1;
wire na1680_2;
wire na1682_1;
wire na1682_4;
wire na1683_1;
wire na1683_2;
wire na1683_4;
wire na1685_1;
wire na1685_2;
wire na1687_1;
wire na1687_4;
wire na1688_1;
wire na1688_2;
wire na1688_4;
wire na1690_1;
wire na1690_2;
wire na1690_4;
wire na1692_1;
wire na1693_1;
wire na1693_4;
wire na1694_1;
wire na1694_2;
wire na1694_4;
wire na1696_1;
wire na1696_2;
wire na1696_4;
wire na1698_1;
wire na1699_4;
wire na1701_1;
wire na1701_4;
wire na1702_4;
wire na1704_1;
wire na1704_4;
wire na1705_1;
wire na1705_2;
wire na1705_4;
wire na1707_1;
wire na1708_1;
wire na1708_4;
wire na1709_1;
wire na1709_2;
wire na1709_4;
wire na1711_1;
wire na1711_2;
wire na1713_1;
wire na1713_4;
wire na1714_1;
wire na1714_2;
wire na1714_4;
wire na1716_1;
wire na1716_2;
wire na1718_1;
wire na1718_2;
wire na1718_4;
wire na1720_1;
wire na1721_1;
wire na1721_4;
wire na1722_1;
wire na1722_2;
wire na1722_4;
wire na1724_1;
wire na1724_2;
wire na1724_4;
wire na1726_1;
wire na1727_1;
wire na1727_4;
wire na1728_1;
wire na1728_2;
wire na1728_4;
wire na1730_1;
wire na1730_2;
wire na1732_1;
wire na1732_4;
wire na1733_1;
wire na1733_2;
wire na1733_4;
wire na1735_1;
wire na1735_2;
wire na1739_1;
wire na1739_2;
wire na1741_1;
wire na1741_1_i;
wire na1741_2;
wire na1741_2_i;
wire na1743_1;
wire na1743_1_i;
wire na1743_2;
wire na1743_2_i;
wire na1745_1;
wire na1745_1_i;
wire na1745_2;
wire na1745_2_i;
wire na1747_1;
wire na1747_1_i;
wire na1747_2;
wire na1747_2_i;
wire na1763_1;
wire na1763_1_i;
wire na1763_2;
wire na1763_2_i;
wire na1765_1;
wire na1765_1_i;
wire na1765_2;
wire na1765_2_i;
wire na1767_1;
wire na1767_1_i;
wire na1767_2;
wire na1767_2_i;
wire na1769_1;
wire na1769_1_i;
wire na1769_2;
wire na1769_2_i;
wire na1771_1;
wire na1771_1_i;
wire na1771_2;
wire na1771_2_i;
wire na1773_1;
wire na1773_1_i;
wire na1773_2;
wire na1773_2_i;
wire na1775_1;
wire na1775_1_i;
wire na1775_2;
wire na1775_2_i;
wire na1777_1;
wire na1777_1_i;
wire na1777_2;
wire na1777_2_i;
wire na1780_1;
wire na1780_1_i;
wire na1780_2;
wire na1780_2_i;
wire na1782_1;
wire na1782_1_i;
wire na1782_2;
wire na1782_2_i;
wire na1784_1;
wire na1784_1_i;
wire na1784_2;
wire na1784_2_i;
wire na1786_1;
wire na1786_1_i;
wire na1786_2;
wire na1786_2_i;
wire na1788_1;
wire na1788_1_i;
wire na1788_2;
wire na1788_2_i;
wire na1790_1;
wire na1790_1_i;
wire na1790_2;
wire na1790_2_i;
wire na1792_1;
wire na1792_1_i;
wire na1792_2;
wire na1792_2_i;
wire na1794_1;
wire na1794_1_i;
wire na1794_2;
wire na1794_2_i;
wire na1811_1;
wire na1811_1_i;
wire na1811_2;
wire na1811_2_i;
wire na1813_1;
wire na1813_1_i;
wire na1813_2;
wire na1813_2_i;
wire na1815_1;
wire na1815_1_i;
wire na1815_2;
wire na1815_2_i;
wire na1817_1;
wire na1817_1_i;
wire na1817_2;
wire na1817_2_i;
wire na1819_1;
wire na1819_1_i;
wire na1819_2;
wire na1819_2_i;
wire na1821_1;
wire na1821_1_i;
wire na1821_2;
wire na1821_2_i;
wire na1823_1;
wire na1823_1_i;
wire na1823_2;
wire na1823_2_i;
wire na1825_1;
wire na1825_1_i;
wire na1825_2;
wire na1825_2_i;
wire na1862_1;
wire na1862_1_i;
wire na1862_2;
wire na1862_2_i;
wire na1864_1;
wire na1864_1_i;
wire na1864_2;
wire na1864_2_i;
wire na1866_1;
wire na1866_1_i;
wire na1866_2;
wire na1866_2_i;
wire na1868_1;
wire na1868_1_i;
wire na1868_2;
wire na1868_2_i;
wire na1878_1;
wire na1878_1_i;
wire na1878_2;
wire na1878_2_i;
wire na1880_1;
wire na1880_1_i;
wire na1880_2;
wire na1880_2_i;
wire na1882_1;
wire na1882_1_i;
wire na1882_2;
wire na1882_2_i;
wire na1884_1;
wire na1884_1_i;
wire na1884_2;
wire na1884_2_i;
wire na1887_1;
wire na1887_1_i;
wire na1887_2;
wire na1887_2_i;
wire na1889_1;
wire na1889_1_i;
wire na1889_2;
wire na1889_2_i;
wire na1891_1;
wire na1891_1_i;
wire na1891_2;
wire na1891_2_i;
wire na1893_1;
wire na1893_1_i;
wire na1893_2;
wire na1893_2_i;
wire na1984_2;
wire na1984_2_i;
wire na1985_1;
wire na1985_1_i;
wire na1986_1;
wire na1986_1_i;
wire na1986_2;
wire na1986_2_i;
wire na1989_2;
wire na1989_2_i;
wire na1990_1;
wire na1990_1_i;
wire na1990_2;
wire na1990_2_i;
wire na1991_1;
wire na1991_1_i;
wire na1993_1;
wire na1993_1_i;
wire na1993_2;
wire na1993_2_i;
wire na1994_2;
wire na1994_2_i;
wire na1995_1;
wire na1995_1_i;
wire na1996_2;
wire na1996_2_i;
wire na1997_1;
wire na1997_1_i;
wire na1998_2;
wire na1998_2_i;
wire na1999_1;
wire na1999_1_i;
wire na2000_2;
wire na2000_2_i;
wire na2001_1;
wire na2001_1_i;
wire na2001_2;
wire na2001_2_i;
wire na2002_1;
wire na2002_1_i;
wire na2011_1;
wire na2011_1_i;
wire na2011_2;
wire na2011_2_i;
wire na2013_1;
wire na2013_1_i;
wire na2013_2;
wire na2013_2_i;
wire na2015_1;
wire na2015_1_i;
wire na2015_2;
wire na2015_2_i;
wire na2017_1;
wire na2017_1_i;
wire na2017_2;
wire na2017_2_i;
wire na2019_1;
wire na2019_1_i;
wire na2019_2;
wire na2019_2_i;
wire na2021_1;
wire na2021_1_i;
wire na2021_2;
wire na2021_2_i;
wire na2023_1;
wire na2023_1_i;
wire na2023_2;
wire na2023_2_i;
wire na2025_1;
wire na2025_1_i;
wire na2025_2;
wire na2025_2_i;
wire na2027_1;
wire na2027_1_i;
wire na2027_2;
wire na2027_2_i;
wire na2029_1;
wire na2029_1_i;
wire na2029_2;
wire na2029_2_i;
wire na2031_1;
wire na2031_1_i;
wire na2031_2;
wire na2031_2_i;
wire na2033_1;
wire na2033_1_i;
wire na2033_2;
wire na2033_2_i;
wire na2035_1;
wire na2035_1_i;
wire na2035_2;
wire na2035_2_i;
wire na2037_1;
wire na2037_1_i;
wire na2037_2;
wire na2037_2_i;
wire na2039_1;
wire na2039_1_i;
wire na2039_2;
wire na2039_2_i;
wire na2041_2;
wire na2041_2_i;
wire na2091_1;
wire na2091_1_i;
wire na2091_2;
wire na2091_2_i;
wire na2093_1;
wire na2093_1_i;
wire na2118_1;
wire na2118_1_i;
wire na2118_2;
wire na2118_2_i;
wire na2120_1;
wire na2120_1_i;
wire na2120_2;
wire na2120_2_i;
wire na2122_1;
wire na2122_1_i;
wire na2122_2;
wire na2122_2_i;
wire na2124_1;
wire na2124_1_i;
wire na2124_2;
wire na2124_2_i;
wire na2125_1;
wire na2125_1_i;
wire na2125_2;
wire na2125_2_i;
wire na2127_1;
wire na2127_1_i;
wire na2127_2;
wire na2127_2_i;
wire na2129_1;
wire na2129_1_i;
wire na2129_2;
wire na2129_2_i;
wire na2221_2;
wire na2221_2_i;
wire na2222_1;
wire na2222_1_i;
wire na2223_1;
wire na2223_1_i;
wire na2223_2;
wire na2223_2_i;
wire na2226_2;
wire na2226_2_i;
wire na2228_1;
wire na2228_1_i;
wire na2228_2;
wire na2228_2_i;
wire na2229_1;
wire na2229_1_i;
wire na2229_2;
wire na2229_2_i;
wire na2230_1;
wire na2230_1_i;
wire na2231_1;
wire na2231_1_i;
wire na2232_1;
wire na2232_1_i;
wire na2233_2;
wire na2233_2_i;
wire na2234_1;
wire na2234_1_i;
wire na2235_2;
wire na2235_2_i;
wire na2236_1;
wire na2236_1_i;
wire na2237_2;
wire na2237_2_i;
wire na2238_1;
wire na2238_1_i;
wire na2238_2;
wire na2238_2_i;
wire na2239_1;
wire na2239_1_i;
wire na2246_2;
wire na2246_2_i;
wire na2248_1;
wire na2248_1_i;
wire na2248_2;
wire na2248_2_i;
wire na2250_1;
wire na2250_1_i;
wire na2250_2;
wire na2250_2_i;
wire na2252_1;
wire na2252_1_i;
wire na2252_2;
wire na2252_2_i;
wire na2254_1;
wire na2254_1_i;
wire na2254_2;
wire na2254_2_i;
wire na2256_1;
wire na2256_1_i;
wire na2256_2;
wire na2256_2_i;
wire na2258_1;
wire na2258_1_i;
wire na2258_2;
wire na2258_2_i;
wire na2260_1;
wire na2260_1_i;
wire na2260_2;
wire na2260_2_i;
wire na2262_1;
wire na2262_1_i;
wire na2262_2;
wire na2262_2_i;
wire na2264_1;
wire na2264_1_i;
wire na2264_2;
wire na2264_2_i;
wire na2266_1;
wire na2266_1_i;
wire na2266_2;
wire na2266_2_i;
wire na2268_1;
wire na2268_1_i;
wire na2268_2;
wire na2268_2_i;
wire na2270_1;
wire na2270_1_i;
wire na2270_2;
wire na2270_2_i;
wire na2272_1;
wire na2272_1_i;
wire na2272_2;
wire na2272_2_i;
wire na2274_1;
wire na2274_1_i;
wire na2274_2;
wire na2274_2_i;
wire na2276_1;
wire na2276_1_i;
wire na2276_2;
wire na2276_2_i;
wire na2278_2;
wire na2278_2_i;
wire na2337_1;
wire na2337_1_i;
wire na2337_2;
wire na2337_2_i;
wire na2339_1;
wire na2339_1_i;
wire na2350_2;
wire na2350_2_i;
wire na2352_1;
wire na2352_1_i;
wire na2352_2;
wire na2352_2_i;
wire na2354_1;
wire na2354_1_i;
wire na2354_2;
wire na2354_2_i;
wire na2356_1;
wire na2356_1_i;
wire na2356_2;
wire na2356_2_i;
wire na2358_1;
wire na2358_1_i;
wire na2358_2;
wire na2358_2_i;
wire na2359_1;
wire na2359_1_i;
wire na2359_2;
wire na2359_2_i;
wire na2361_1;
wire na2361_1_i;
wire na2361_2;
wire na2361_2_i;
wire na2363_1;
wire na2363_1_i;
wire na2363_2;
wire na2363_2_i;
wire na2472_1;
wire na2472_1_i;
wire na2473_2;
wire na2473_2_i;
wire na2474_1;
wire na2474_1_i;
wire na2474_2;
wire na2474_2_i;
wire na2477_1;
wire na2477_1_i;
wire na2478_1;
wire na2478_1_i;
wire na2478_2;
wire na2478_2_i;
wire na2479_2;
wire na2479_2_i;
wire na2481_1;
wire na2481_1_i;
wire na2481_2;
wire na2481_2_i;
wire na2482_1;
wire na2482_1_i;
wire na2483_2;
wire na2483_2_i;
wire na2484_1;
wire na2484_1_i;
wire na2485_2;
wire na2485_2_i;
wire na2486_1;
wire na2486_1_i;
wire na2487_2;
wire na2487_2_i;
wire na2488_1;
wire na2488_1_i;
wire na2489_1;
wire na2489_1_i;
wire na2489_2;
wire na2489_2_i;
wire na2490_2;
wire na2490_2_i;
wire na2497_1;
wire na2497_1_i;
wire na2499_1;
wire na2499_1_i;
wire na2499_2;
wire na2499_2_i;
wire na2501_1;
wire na2501_1_i;
wire na2501_2;
wire na2501_2_i;
wire na2503_1;
wire na2503_1_i;
wire na2503_2;
wire na2503_2_i;
wire na2505_1;
wire na2505_1_i;
wire na2505_2;
wire na2505_2_i;
wire na2507_1;
wire na2507_1_i;
wire na2507_2;
wire na2507_2_i;
wire na2509_1;
wire na2509_1_i;
wire na2509_2;
wire na2509_2_i;
wire na2511_1;
wire na2511_1_i;
wire na2511_2;
wire na2511_2_i;
wire na2513_1;
wire na2513_1_i;
wire na2513_2;
wire na2513_2_i;
wire na2515_1;
wire na2515_1_i;
wire na2515_2;
wire na2515_2_i;
wire na2517_1;
wire na2517_1_i;
wire na2517_2;
wire na2517_2_i;
wire na2519_1;
wire na2519_1_i;
wire na2519_2;
wire na2519_2_i;
wire na2521_1;
wire na2521_1_i;
wire na2521_2;
wire na2521_2_i;
wire na2523_1;
wire na2523_1_i;
wire na2523_2;
wire na2523_2_i;
wire na2525_1;
wire na2525_1_i;
wire na2525_2;
wire na2525_2_i;
wire na2527_1;
wire na2527_1_i;
wire na2527_2;
wire na2527_2_i;
wire na2529_2;
wire na2529_2_i;
wire na2579_1;
wire na2579_1_i;
wire na2579_2;
wire na2579_2_i;
wire na2581_1;
wire na2581_1_i;
wire na2593_1;
wire na2593_1_i;
wire na2593_2;
wire na2593_2_i;
wire na2595_1;
wire na2595_1_i;
wire na2595_2;
wire na2595_2_i;
wire na2597_1;
wire na2597_1_i;
wire na2597_2;
wire na2597_2_i;
wire na2599_1;
wire na2599_1_i;
wire na2599_2;
wire na2599_2_i;
wire na2600_1;
wire na2600_1_i;
wire na2600_2;
wire na2600_2_i;
wire na2602_1;
wire na2602_1_i;
wire na2602_2;
wire na2602_2_i;
wire na2604_1;
wire na2604_1_i;
wire na2604_2;
wire na2604_2_i;
wire na2705_2;
wire na2705_2_i;
wire na2706_1;
wire na2706_1_i;
wire na2707_1;
wire na2707_1_i;
wire na2707_2;
wire na2707_2_i;
wire na2710_2;
wire na2710_2_i;
wire na2712_1;
wire na2712_1_i;
wire na2712_2;
wire na2712_2_i;
wire na2713_1;
wire na2713_1_i;
wire na2713_2;
wire na2713_2_i;
wire na2714_1;
wire na2714_1_i;
wire na2715_2;
wire na2715_2_i;
wire na2716_1;
wire na2716_1_i;
wire na2717_2;
wire na2717_2_i;
wire na2718_1;
wire na2718_1_i;
wire na2719_2;
wire na2719_2_i;
wire na2720_1;
wire na2720_1_i;
wire na2721_2;
wire na2721_2_i;
wire na2722_1;
wire na2722_1_i;
wire na2722_2;
wire na2722_2_i;
wire na2723_2;
wire na2723_2_i;
wire na2730_2;
wire na2730_2_i;
wire na2739_1;
wire na2739_1_i;
wire na2739_2;
wire na2739_2_i;
wire na2741_1;
wire na2741_1_i;
wire na2741_2;
wire na2741_2_i;
wire na2743_1;
wire na2743_1_i;
wire na2743_2;
wire na2743_2_i;
wire na2745_1;
wire na2745_1_i;
wire na2745_2;
wire na2745_2_i;
wire na2747_1;
wire na2747_1_i;
wire na2747_2;
wire na2747_2_i;
wire na2749_1;
wire na2749_1_i;
wire na2749_2;
wire na2749_2_i;
wire na2751_1;
wire na2751_1_i;
wire na2751_2;
wire na2751_2_i;
wire na2753_1;
wire na2753_1_i;
wire na2753_2;
wire na2753_2_i;
wire na2755_1;
wire na2755_1_i;
wire na2755_2;
wire na2755_2_i;
wire na2757_1;
wire na2757_1_i;
wire na2757_2;
wire na2757_2_i;
wire na2759_1;
wire na2759_1_i;
wire na2759_2;
wire na2759_2_i;
wire na2761_1;
wire na2761_1_i;
wire na2761_2;
wire na2761_2_i;
wire na2763_1;
wire na2763_1_i;
wire na2763_2;
wire na2763_2_i;
wire na2765_1;
wire na2765_1_i;
wire na2765_2;
wire na2765_2_i;
wire na2767_1;
wire na2767_1_i;
wire na2767_2;
wire na2767_2_i;
wire na2769_1;
wire na2769_1_i;
wire na2819_1;
wire na2819_1_i;
wire na2819_2;
wire na2819_2_i;
wire na2821_2;
wire na2821_2_i;
wire na2840_1;
wire na2840_1_i;
wire na2840_2;
wire na2840_2_i;
wire na2842_1;
wire na2842_1_i;
wire na2842_2;
wire na2842_2_i;
wire na2844_1;
wire na2844_1_i;
wire na2844_2;
wire na2844_2_i;
wire na2846_1;
wire na2846_1_i;
wire na2846_2;
wire na2846_2_i;
wire na2847_1;
wire na2847_1_i;
wire na2847_2;
wire na2847_2_i;
wire na2849_1;
wire na2849_1_i;
wire na2849_2;
wire na2849_2_i;
wire na2851_1;
wire na2851_1_i;
wire na2851_2;
wire na2851_2_i;
wire na2956_1;
wire na2956_1_i;
wire na2957_2;
wire na2957_2_i;
wire na2958_1;
wire na2958_1_i;
wire na2958_2;
wire na2958_2_i;
wire na2961_1;
wire na2961_1_i;
wire na2962_1;
wire na2962_1_i;
wire na2962_2;
wire na2962_2_i;
wire na2963_2;
wire na2963_2_i;
wire na2965_1;
wire na2965_1_i;
wire na2965_2;
wire na2965_2_i;
wire na2966_1;
wire na2966_1_i;
wire na2967_2;
wire na2967_2_i;
wire na2968_1;
wire na2968_1_i;
wire na2969_2;
wire na2969_2_i;
wire na2970_1;
wire na2970_1_i;
wire na2971_2;
wire na2971_2_i;
wire na2972_1;
wire na2972_1_i;
wire na2973_1;
wire na2973_1_i;
wire na2973_2;
wire na2973_2_i;
wire na2974_2;
wire na2974_2_i;
wire na2981_1;
wire na2981_1_i;
wire na2984_1;
wire na2984_1_i;
wire na2984_2;
wire na2984_2_i;
wire na2986_1;
wire na2986_1_i;
wire na2986_2;
wire na2986_2_i;
wire na2988_1;
wire na2988_1_i;
wire na2988_2;
wire na2988_2_i;
wire na2990_1;
wire na2990_1_i;
wire na2990_2;
wire na2990_2_i;
wire na2992_1;
wire na2992_1_i;
wire na2992_2;
wire na2992_2_i;
wire na2994_1;
wire na2994_1_i;
wire na2994_2;
wire na2994_2_i;
wire na2996_1;
wire na2996_1_i;
wire na2996_2;
wire na2996_2_i;
wire na2998_1;
wire na2998_1_i;
wire na2998_2;
wire na2998_2_i;
wire na3000_1;
wire na3000_1_i;
wire na3000_2;
wire na3000_2_i;
wire na3002_1;
wire na3002_1_i;
wire na3002_2;
wire na3002_2_i;
wire na3004_1;
wire na3004_1_i;
wire na3004_2;
wire na3004_2_i;
wire na3006_1;
wire na3006_1_i;
wire na3006_2;
wire na3006_2_i;
wire na3008_1;
wire na3008_1_i;
wire na3008_2;
wire na3008_2_i;
wire na3010_1;
wire na3010_1_i;
wire na3010_2;
wire na3010_2_i;
wire na3012_1;
wire na3012_1_i;
wire na3012_2;
wire na3012_2_i;
wire na3014_2;
wire na3014_2_i;
wire na3064_1;
wire na3064_1_i;
wire na3064_2;
wire na3064_2_i;
wire na3066_1;
wire na3066_1_i;
wire na3098_1;
wire na3098_1_i;
wire na3098_2;
wire na3098_2_i;
wire na3100_1;
wire na3100_1_i;
wire na3100_2;
wire na3100_2_i;
wire na3102_1;
wire na3102_1_i;
wire na3102_2;
wire na3102_2_i;
wire na3104_1;
wire na3104_1_i;
wire na3104_2;
wire na3104_2_i;
wire na3105_1;
wire na3105_1_i;
wire na3105_2;
wire na3105_2_i;
wire na3107_1;
wire na3107_1_i;
wire na3107_2;
wire na3107_2_i;
wire na3109_1;
wire na3109_1_i;
wire na3109_2;
wire na3109_2_i;
wire na3145_1;
wire na3146_1;
wire na3147_1;
wire na3148_1;
wire na3149_1;
wire na3150_1;
wire na3151_1;
wire na3152_1;
wire na3153_1;
wire na3154_1;
wire na3155_1;
wire na3156_1;
wire na3157_1;
wire na3158_1;
wire na3159_1;
wire na3160_1;
wire na3161_1;
wire na3162_1;
wire na3163_2;
wire na3164_1;
wire na3165_1;
wire na3166_1;
wire na3167_1;
wire na3168_1;
wire na3169_1;
wire na3170_1;
wire na3171_1;
wire na3172_1;
wire na3173_1;
wire na3174_1;
wire na3175_1;
wire na3176_1;
wire na3177_1;
wire na3178_1;
wire na3179_1;
wire na3180_1;
wire na3181_1;
wire na3182_1;
wire na3183_1;
wire na3184_1;
wire na3185_1;
wire na3186_1;
wire na3187_1;
wire na3188_1;
wire na3189_1;
wire na3190_1;
wire na3191_1;
wire na3192_1;
wire na3193_1;
wire na3194_1;
wire na3195_1;
wire na3196_1;
wire na3197_1;
wire na3198_1;
wire na3199_1;
wire na3200_1;
wire na3201_1;
wire na3202_1;
wire na3203_1;
wire na3204_1;
wire na3205_1;
wire na3206_1;
wire na3207_1;
wire na3208_1;
wire na3209_1;
wire na3210_1;
wire na3211_1;
wire na3212_1;
wire na3213_1;
wire na3214_1;
wire na3215_1;
wire na3216_1;
wire na3217_1;
wire na3218_1;
wire na3219_1;
wire na3220_1;
wire na3222_2;
wire na3222_3;
wire na3222_4;
wire na3222_5;
wire na3222_6;
wire na3224_2;
wire na3227_2;
wire na3228_1;
wire na3229_1;
wire na3229_2;
wire na3230_2;
wire na3231_2;
wire na3232_2;
wire na3233_1;
wire na3233_9;
wire na3234_1;
wire na3234_4;
wire na3235_1;
wire na3235_4;
wire na3236_2;
wire na3237_1;
wire na3237_9;
wire na3238_2;
wire na3239_1;
wire na3239_9;
wire na3240_2;
wire na3241_2;
wire na3242_1;
wire na3242_9;
wire na3243_1;
wire na3244_2;
wire na3245_1;
wire na3245_9;
wire na3246_1;
wire na3247_1;
wire na3247_4;
wire na3248_1;
wire na3249_1;
wire na3250_2;
wire na3251_1;
wire na3251_9;
wire na3252_1;
wire na3253_2;
wire na3254_2;
wire na3255_1;
wire na3256_2;
wire na3257_1;
wire na3257_9;
wire na3258_1;
wire na3258_2;
wire na3259_1;
wire na3260_1;
wire na3260_4;
wire na3261_2;
wire na3262_1;
wire na3263_1;
wire na3264_1;
wire na3264_9;
wire na3265_2;
wire na3266_1;
wire na3266_9;
wire na3267_1;
wire na3267_4;
wire na3268_1;
wire na3268_2;
wire na3269_2;
wire na3270_2;
wire na3271_1;
wire na3271_9;
wire na3272_1;
wire na3273_2;
wire na3274_2;
wire na3275_1;
wire na3276_1;
wire na3277_1;
wire na3277_9;
wire na3278_1;
wire na3278_2;
wire na3279_1;
wire na3280_2;
wire na3281_1;
wire na3281_4;
wire na3282_1;
wire na3283_1;
wire na3284_1;
wire na3284_9;
wire na3285_1;
wire na3286_2;
wire na3287_1;
wire na3288_1;
wire na3289_1;
wire na3289_9;
wire na3290_1;
wire na3290_2;
wire na3291_2;
wire na3292_1;
wire na3293_1;
wire na3293_9;
wire na3294_2;
wire na3295_1;
wire na3295_9;
wire na3296_1;
wire na3296_2;
wire na3297_2;
wire na3298_1;
wire na3299_1;
wire na3299_9;
wire na3300_2;
wire na3301_1;
wire na3302_2;
wire na3303_1;
wire na3304_1;
wire na3304_9;
wire na3305_2;
wire na3306_2;
wire na3307_2;
wire na3308_1;
wire na3308_9;
wire na3309_2;
wire na3310_1;
wire na3311_1;
wire na3311_9;
wire na3312_1;
wire na3313_1;
wire na3314_2;
wire na3315_1;
wire na3315_9;
wire na3316_1;
wire na3317_1;
wire na3318_2;
wire na3319_1;
wire na3319_9;
wire na3320_2;
wire na3321_1;
wire na3321_9;
wire na3322_1;
wire na3322_2;
wire na3323_2;
wire na3324_1;
wire na3325_1;
wire na3325_9;
wire na3326_2;
wire na3327_1;
wire na3328_2;
wire na3329_2;
wire na3330_1;
wire na3330_9;
wire na3331_1;
wire na3332_2;
wire na3333_1;
wire na3333_9;
wire na3334_1;
wire na3335_1;
wire na3336_1;
wire na3337_2;
wire na3338_2;
wire na3339_1;
wire na3339_9;
wire na3340_2;
wire na3341_1;
wire na3342_2;
wire na3343_1;
wire na3344_1;
wire na3344_9;
wire na3345_2;
wire na3346_1;
wire na3347_1;
wire na3347_9;
wire na3348_1;
wire na3349_2;
wire na3350_1;
wire na3350_9;
wire na3351_2;
wire na3352_1;
wire na3352_9;
wire na3353_2;
wire na3354_1;
wire na3354_9;
wire na3355_2;
wire na3356_1;
wire na3356_9;
wire na3357_2;
wire na3358_1;
wire na3358_9;
wire na3359_2;
wire na3360_1;
wire na3360_9;
wire na3361_2;
wire na3362_1;
wire na3362_9;
wire na3363_2;
wire na3364_1;
wire na3364_9;
wire na3365_2;
wire na3366_1;
wire na3366_9;
wire na3367_2;
wire na3368_1;
wire na3368_9;
wire na3369_2;
wire na3370_1;
wire na3370_9;
wire na3371_2;
wire na3372_1;
wire na3372_9;
wire na3373_2;
wire na3374_1;
wire na3374_9;
wire na3375_2;
wire na3376_1;
wire na3376_9;
wire na3377_2;
wire na3378_1;
wire na3378_9;
wire na3379_2;
wire na3380_1;
wire na3380_9;
wire na3381_2;
wire na3382_1;
wire na3382_9;
wire na3383_2;
wire na3384_1;
wire na3384_9;
wire na3385_2;
wire na3386_1;
wire na3386_9;
wire na3387_2;
wire na3388_1;
wire na3388_9;
wire na3389_2;
wire na3390_1;
wire na3390_9;
wire na3391_2;
wire na3392_1;
wire na3392_9;
wire na3393_2;
wire na3394_1;
wire na3394_9;
wire na3395_2;
wire na3396_1;
wire na3396_9;
wire na3397_2;
wire na3398_1;
wire na3398_9;
wire na3399_2;
wire na3400_1;
wire na3400_9;
wire na3401_2;
wire na3402_1;
wire na3402_9;
wire na3403_2;
wire na3404_1;
wire na3404_9;
wire na3405_2;
wire na3406_1;
wire na3406_9;
wire na3407_2;
wire na3408_1;
wire na3408_9;
wire na3409_2;
wire na3410_1;
wire na3410_9;
wire na3411_2;
wire na3412_1;
wire na3412_9;
wire na3413_2;
wire na3414_1;
wire na3415_1;
wire na3416_2;
wire na3417_1;
wire na3418_1;
wire na3419_1;
wire na3420_2;
wire na3421_1;
wire na3422_1;
wire na3423_2;
wire na3424_1;
wire na3425_1;
wire na3426_2;
wire na3427_1;
wire na3428_1;
wire na3429_2;
wire na3430_1;
wire na3431_1;
wire na3432_1;
wire na3433_2;
wire na3434_2;
wire na3435_2;
wire na3436_1;
wire na3437_1;
wire na3438_1;
wire na3439_2;
wire na3440_1;
wire na3441_2;
wire na3442_1;
wire na3443_2;
wire na3444_1;
wire na3445_2;
wire na3446_2;
wire na3447_2;
wire na3448_1;
wire na3449_2;
wire na3450_1;
wire na3450_9;
wire na3451_1;
wire na3451_2;
wire na3452_2;
wire na3453_1;
wire na3453_2;
wire na3454_2;
wire na3455_1;
wire na3455_9;
wire na3456_2;
wire na3457_1;
wire na3458_2;
wire na3459_1;
wire na3460_1;
wire na3460_9;
wire na3461_1;
wire na3462_1;
wire na3463_1;
wire na3464_1;
wire na3465_1;
wire na3466_2;
wire na3467_2;
wire na3468_2;
wire na3469_1;
wire na3469_9;
wire na3470_1;
wire na3471_2;
wire na3472_1;
wire na3473_2;
wire na3474_1;
wire na3474_9;
wire na3475_2;
wire na3476_1;
wire na3476_9;
wire na3477_2;
wire na3478_1;
wire na3478_9;
wire na3479_2;
wire na3480_1;
wire na3480_9;
wire na3481_2;
wire na3482_1;
wire na3482_9;
wire na3483_2;
wire na3484_1;
wire na3484_9;
wire na3485_2;
wire na3486_1;
wire na3486_9;
wire na3487_2;
wire na3488_1;
wire na3488_9;
wire na3489_2;
wire na3490_1;
wire na3490_9;
wire na3491_2;
wire na3492_1;
wire na3492_9;
wire na3493_2;
wire na3494_1;
wire na3494_9;
wire na3495_2;
wire na3496_1;
wire na3496_9;
wire na3497_2;
wire na3498_1;
wire na3498_9;
wire na3499_2;
wire na3500_1;
wire na3500_9;
wire na3501_2;
wire na3502_1;
wire na3502_9;
wire na3503_2;
wire na3504_1;
wire na3504_9;
wire na3505_2;
wire na3506_1;
wire na3506_9;
wire na3507_2;
wire na3508_1;
wire na3508_9;
wire na3509_2;
wire na3510_1;
wire na3510_9;
wire na3511_2;
wire na3512_1;
wire na3512_9;
wire na3513_2;
wire na3514_1;
wire na3514_9;
wire na3515_2;
wire na3516_1;
wire na3516_9;
wire na3517_2;
wire na3518_1;
wire na3518_9;
wire na3519_2;
wire na3520_1;
wire na3520_9;
wire na3521_2;
wire na3522_1;
wire na3522_9;
wire na3523_2;
wire na3524_1;
wire na3524_9;
wire na3525_2;
wire na3526_1;
wire na3527_2;
wire na3528_1;
wire na3529_2;
wire na3530_1;
wire na3531_2;
wire na3532_1;
wire na3533_2;
wire na3534_2;
wire na3535_2;
wire na3536_1;
wire na3536_9;
wire na3537_2;
wire na3538_1;
wire na3538_9;
wire na3539_1;
wire na3540_2;
wire na3541_1;
wire na3541_9;
wire na3542_1;
wire na3543_1;
wire na3544_2;
wire na3545_1;
wire na3545_9;
wire na3546_1;
wire na3547_2;
wire na3548_1;
wire na3548_9;
wire na3549_1;
wire na3550_2;
wire na3551_1;
wire na3551_9;
wire na3552_1;
wire na3553_2;
wire na3554_1;
wire na3554_9;
wire na3555_1;
wire na3556_2;
wire na3557_2;
wire na3558_2;
wire na3559_1;
wire na3560_1;
wire na3561_1;
wire na3562_2;
wire na3563_2;
wire na3564_1;
wire na3565_2;
wire na3566_1;
wire na3566_9;
wire na3567_2;
wire na3568_1;
wire na3568_9;
wire na3569_2;
wire na3570_2;
wire na3571_1;
wire na3571_2;
wire na3572_1;
wire na3572_9;
wire na3573_2;
wire na3574_1;
wire na3574_9;
wire na3575_1;
wire na3576_2;
wire na3577_2;
wire na3578_1;
wire na3579_1;
wire na3579_9;
wire na3580_1;
wire na3581_2;
wire na3582_1;
wire na3583_1;
wire na3583_9;
wire na3584_2;
wire na3585_1;
wire na3586_1;
wire na3586_9;
wire na3587_2;
wire na3588_1;
wire na3589_1;
wire na3590_1;
wire na3591_1;
wire na3591_9;
wire na3592_2;
wire na3593_1;
wire na3593_9;
wire na3594_2;
wire na3595_1;
wire na3595_9;
wire na3596_2;
wire na3597_1;
wire na3597_9;
wire na3598_2;
wire na3599_1;
wire na3599_9;
wire na3600_2;
wire na3601_1;
wire na3601_9;
wire na3602_2;
wire na3603_1;
wire na3603_9;
wire na3604_2;
wire na3605_1;
wire na3605_9;
wire na3606_2;
wire na3607_1;
wire na3607_9;
wire na3608_2;
wire na3609_1;
wire na3609_9;
wire na3610_2;
wire na3611_1;
wire na3611_9;
wire na3612_2;
wire na3613_1;
wire na3613_9;
wire na3614_2;
wire na3615_1;
wire na3615_9;
wire na3616_2;
wire na3617_1;
wire na3617_9;
wire na3618_2;
wire na3619_1;
wire na3619_9;
wire na3620_2;
wire na3621_1;
wire na3621_9;
wire na3622_2;
wire na3623_1;
wire na3623_9;
wire na3624_2;
wire na3625_1;
wire na3625_9;
wire na3626_2;
wire na3627_1;
wire na3627_9;
wire na3628_2;
wire na3629_1;
wire na3629_9;
wire na3630_2;
wire na3631_1;
wire na3631_9;
wire na3632_2;
wire na3633_1;
wire na3633_9;
wire na3634_2;
wire na3635_1;
wire na3635_9;
wire na3636_2;
wire na3637_1;
wire na3637_9;
wire na3638_2;
wire na3639_1;
wire na3639_9;
wire na3640_2;
wire na3641_1;
wire na3641_9;
wire na3642_2;
wire na3643_1;
wire na3643_9;
wire na3644_2;
wire na3645_1;
wire na3645_9;
wire na3646_2;
wire na3647_1;
wire na3647_9;
wire na3648_2;
wire na3649_1;
wire na3649_9;
wire na3650_2;
wire na3651_1;
wire na3651_9;
wire na3652_2;
wire na3653_1;
wire na3653_9;
wire na3654_2;
wire na3655_1;
wire na3655_9;
wire na3656_2;
wire na3657_2;
wire na3658_1;
wire na3658_9;
wire na3659_2;
wire na3660_2;
wire na3661_1;
wire na3662_1;
wire na3662_9;
wire na3663_2;
wire na3664_1;
wire na3665_1;
wire na3665_9;
wire na3666_2;
wire na3667_1;
wire na3668_1;
wire na3668_9;
wire na3669_2;
wire na3670_1;
wire na3671_1;
wire na3671_9;
wire na3672_2;
wire na3673_1;
wire na3674_2;
wire na3675_1;
wire na3676_1;
wire na3677_1;
wire na3678_2;
wire na3679_1;
wire na3680_1;
wire na3681_1;
wire na3681_9;
wire na3682_1;
wire na3683_1;
wire na3684_2;
wire na3685_1;
wire na3685_9;
wire na3686_2;
wire na3687_1;
wire na3687_9;
wire na3688_2;
wire na3689_1;
wire na3689_2;
wire na3690_2;
wire na3691_1;
wire na3691_9;
wire na3692_2;
wire na3693_1;
wire na3694_2;
wire na3695_1;
wire na3696_1;
wire na3696_9;
wire na3697_2;
wire na3698_1;
wire na3699_2;
wire na3700_1;
wire na3701_2;
wire na3702_1;
wire na3702_9;
wire na3703_1;
wire na3704_2;
wire na3705_1;
wire na3705_9;
wire na3706_1;
wire na3707_1;
wire na3708_2;
wire na3709_2;
wire na3710_1;
wire na3710_9;
wire na3711_2;
wire na3712_1;
wire na3713_2;
wire na3714_1;
wire na3715_2;
wire na3716_1;
wire na3717_2;
wire na3718_1;
wire na3719_2;
wire na3720_1;
wire na3721_2;
wire na3722_1;
wire na3723_2;
wire na3724_1;
wire na3725_2;
wire na3726_1;
wire na3775_2;
wire na3777_2;
wire na3778_1;
wire na3782_1;
wire na3783_1;
wire na3786_1;
wire na3789_1;
wire na3792_1;
wire na3795_1;
wire na3796_1;
wire na3797_2;
wire na3798_2;
wire na3799_2;
wire na3800_1;
wire na3801_1;
wire na3802_1;
wire na3804_1;
wire na3805_2;
wire na3809_1;
wire na3811_2;
wire na3812_1;
wire na3815_1;
wire na3815_2;
wire na3816_2;
wire na3817_1;
wire na3817_2;
wire na3821_1;
wire na3822_2;
wire na3823_1;
wire na3826_1;
wire na3827_1;
wire na3828_1;
wire na3895_1;
wire na3898_2;
wire na3899_1;
wire na3902_1;
wire na3905_1;
wire na3908_1;
wire na3911_1;
wire na3912_2;
wire na3913_2;
wire na3914_1;
wire na3915_1;
wire na3916_1;
wire na3917_2;
wire na3918_2;
wire na3920_1;
wire na3921_2;
wire na3925_1;
wire na3927_2;
wire na3928_1;
wire na3931_1;
wire na3931_2;
wire na3932_1;
wire na3933_1;
wire na3933_2;
wire na3937_1;
wire na3938_1;
wire na3939_1;
wire na3940_2;
wire na3943_1;
wire na3943_2;
wire na3944_2;
wire na3948_1;
wire na3950_2;
wire na3954_1;
wire na3955_2;
wire na3958_1;
wire na3960_2;
wire na3961_2;
wire na3964_1;
wire na3975_1;
wire na3977_1;
wire na3978_1;
wire na3979_1;
wire na3981_1;
wire na3983_1;
wire na3988_1;
wire na3990_1;
wire na3991_1;
wire na3992_1;
wire na3994_1;
wire na3996_2;
wire na4001_1;
wire na4003_1;
wire na4004_1;
wire na4005_1;
wire na4007_1;
wire na4009_1;
wire na4014_1;
wire na4016_1;
wire na4017_1;
wire na4018_1;
wire na4020_1;
wire na4022_2;
wire na4027_1;
wire na4029_1;
wire na4030_1;
wire na4031_1;
wire na4033_1;
wire na4035_2;
wire na4039_1;
wire na4039_2;
wire na4040_1;
wire na4041_1;
wire na4042_2;
wire na4043_1;
wire na4045_1;
wire na4045_2;
wire na4046_1;
wire na4050_1;
wire na4050_2;
wire na4053_1;
wire na4053_2;
wire na4054_2;
wire na4058_1;
wire na4058_2;
wire na4059_2;
wire na4063_1;
wire na4063_2;
wire na4064_1;
wire na4065_2;
wire na4066_2;
wire na4067_2;
wire na4068_2;
wire na4069_2;
wire na4070_2;
wire na4071_2;
wire na4072_2;
wire na4073_2;
wire na4074_2;
wire na4075_2;
wire na4076_2;
wire na4077_2;
wire na4078_2;
wire na4079_2;
wire na4080_2;
wire na4081_2;
wire na4082_2;
wire na4083_2;
wire na4084_2;
wire na4085_2;
wire na4086_2;
wire na4087_2;
wire na4088_2;
wire na4089_2;
wire na4090_2;
wire na4091_2;
wire na4092_2;
wire na4093_2;
wire na4094_2;
wire na4095_2;
wire na4096_2;
wire na4097_2;
wire na4098_2;
wire na4099_2;
wire na4100_2;
wire na4101_2;
wire na4102_2;
wire na4103_2;
wire na4104_2;
wire na4105_2;
wire na4106_2;
wire na4107_2;
wire na4108_2;
wire na4109_2;
wire na4110_2;
wire na4111_2;
wire na4112_2;
wire na4113_2;
wire na4114_2;
wire na4115_2;
wire na4116_2;
wire na4117_2;
wire na4118_2;
wire na4119_2;
wire na4120_2;
wire na4121_2;
wire na4122_2;
wire na4123_2;
wire na4124_2;
wire na4125_2;
wire na4126_2;
wire na4127_2;
wire na4128_2;
wire na4129_2;
wire na4130_2;
wire na4131_2;
wire na4132_2;
wire na4133_2;
wire na4134_2;
wire na4135_2;
wire na4136_2;
wire na4137_2;
wire na4138_2;
wire na4139_2;
wire na4140_2;
wire na4141_2;
wire na4142_2;
wire na4143_2;
wire na4144_2;
wire na4145_2;
wire na4146_2;
wire na4147_2;
wire na4148_2;
wire na4149_2;
wire na4150_2;
wire na4151_2;
wire na4152_2;
wire na4153_2;
wire na4154_2;
wire na4155_2;
wire na4156_2;
wire na4157_2;
wire na4158_2;
wire na4159_2;
wire na4160_2;
wire na4161_2;
wire na4162_2;
wire na4163_2;
wire na4164_2;
wire na4165_2;
wire na4166_2;
wire na4167_2;
wire na4168_2;
wire na4169_2;
wire na4170_2;
wire na4171_2;
wire na4172_2;
wire na4173_2;
wire na4174_2;
wire na4175_2;
wire na4176_2;
wire na4177_2;
wire na4178_2;
wire na4179_2;
wire na4180_2;
wire na4181_2;
wire na4182_2;
wire na4183_2;
wire na4184_2;
wire na4185_2;
wire na4186_2;
wire na4187_2;
wire na4188_2;
wire na4189_2;
wire na4190_2;
wire na4191_2;
wire na4192_2;
wire na4193_2;
wire na4194_2;
wire na4195_2;
wire na4196_2;
wire na4197_2;
wire na4198_2;
wire na4199_2;
wire na4200_2;
wire na4201_2;
wire na4202_2;
wire na4203_2;
wire na4204_2;
wire na4205_2;
wire na4206_2;
wire na4207_2;
wire na4208_2;
wire na4209_2;
wire na4210_2;
wire na4211_2;
wire na4212_2;
wire na4213_2;
wire na4214_2;
wire na4215_2;
wire na4216_2;
wire na4217_2;
wire na4218_2;
wire na4219_2;
wire na4220_2;
wire na4221_2;
wire na4222_2;
wire na4223_2;
wire na4224_2;
wire na4225_2;
wire na4226_2;
wire na4227_2;
wire na4228_2;
wire na4229_2;
wire na4230_2;
wire na4231_2;
wire na4232_2;
wire na4233_2;
wire na4234_2;
wire na4235_2;
wire na4236_2;
wire na4237_2;
wire na4238_2;
wire na4239_2;
wire na4240_2;
wire na4241_2;
wire na4242_2;
wire na4243_2;
wire na4244_2;
wire na4245_2;
wire na4246_2;
wire na4247_2;
wire na4248_2;
wire na4249_2;
wire na4250_2;
wire na4251_2;
wire na4252_2;
wire na4253_2;
wire na4254_2;
wire na4255_2;
wire na4256_2;
wire na4257_2;
wire na4258_2;
wire na4259_2;
wire na4260_2;
wire na4261_2;
wire na4262_2;
wire na4263_2;
wire na4264_2;
wire na4265_2;
wire na4266_2;
wire na4267_2;
wire na4268_2;
wire na4269_2;
wire na4270_2;
wire na4271_2;
wire na4272_2;
wire na4273_2;
wire na4274_2;
wire na4275_2;
wire na4276_2;
wire na4277_2;
wire na4278_2;
wire na4279_2;
wire na4280_2;
wire na4281_2;
wire na4282_2;
wire na4283_2;
wire na4284_2;
wire na4285_2;
wire na4286_2;
wire na4287_2;
wire na4288_2;
wire na4289_2;
wire na4290_2;
wire na4291_2;
wire na4292_2;
wire na4293_2;
wire na4294_2;
wire na4295_2;
wire na4296_2;
wire na4297_2;
wire na4298_2;
wire na4299_2;
wire na4300_2;
wire na4301_2;
wire na4302_2;
wire na4303_2;
wire na4304_2;
wire na4305_2;
wire na4306_2;
wire na4307_2;
wire na4308_2;
wire na4309_2;
wire na4310_2;
wire na4311_2;
wire na4312_2;
wire na4313_2;
wire na4314_2;
wire na4315_2;
wire na4316_2;
wire na4317_2;
wire na4318_2;
wire na4319_2;
wire na4320_2;
wire na4321_2;
wire na4322_2;
wire na4323_2;
wire na4324_2;
wire na4325_2;
wire na4326_2;
wire na4327_2;
wire na4328_2;
wire na4329_2;
wire na4330_2;
wire na4331_2;
wire na4332_2;
wire na4333_2;
wire na4334_2;
wire na4335_2;
wire na4336_2;
wire na4337_2;
wire na4338_2;
wire na4339_2;
wire na4340_2;
wire na4341_2;
wire na4342_2;
wire na4343_2;
wire na4344_2;
wire na4345_2;
wire na4346_2;
wire na4347_2;
wire na4348_2;
wire na4349_2;
wire na4350_2;
wire na4351_2;
wire na4352_2;
wire na4353_2;
wire na4354_2;
wire na4355_2;
wire na4356_2;
wire na4357_2;
wire na4358_2;
wire na4359_2;
wire na4360_2;
wire na4361_2;
wire na4362_2;
wire na4363_2;
wire na4364_2;
wire na4365_2;
wire na4366_2;
wire na4367_2;
wire na4368_2;
wire na4369_2;
wire na4370_2;
wire na4371_2;
wire na4372_2;
wire na4373_2;
wire na4374_2;
wire na4375_2;
wire na4376_2;
wire na4377_2;
wire na4378_2;
wire na4379_2;
wire na4380_2;
wire na4381_2;
wire na4382_2;
wire na4383_2;
wire na4384_2;
wire na4385_2;
wire na4386_2;
wire na4387_2;
wire na4388_2;
wire na4389_2;
wire na4390_2;
wire na4391_2;
wire na4392_2;
wire na4393_2;
wire na4394_2;
wire na4395_2;
wire na4396_2;
wire na4397_2;
wire na4398_2;
wire na4399_2;
wire na4400_2;
wire na4401_2;
wire na4402_2;
wire na4403_2;
wire na4404_2;
wire na4405_2;
wire na4406_2;
wire na4407_2;
wire na4408_2;
wire na4409_2;
wire na4410_2;
wire na4411_2;
wire na4412_2;
wire na4413_2;
wire na4414_2;
wire na4415_2;
wire na4416_2;
wire na4417_2;
wire na4418_2;
wire na4419_2;
wire na4420_2;
wire na4421_2;
wire na4422_2;
wire na4423_2;
wire na4424_2;
wire na4425_2;
wire na4426_2;
wire na4427_2;
wire na4428_2;
wire na4429_2;
wire na4430_2;
wire na4431_2;
wire na4432_2;
wire na4433_2;
wire na4434_2;
wire na4435_2;
wire na4436_2;
wire na4437_2;
wire na4438_2;
wire na4439_2;
wire na4440_2;
wire na4441_2;
wire na4442_2;
wire na4443_2;
wire na4444_2;
wire na4445_2;
wire na4446_2;
wire na4447_2;
wire na4448_2;
wire na4449_2;
wire na4450_2;
wire na4451_2;
wire na4452_2;
wire na4453_2;
wire na4454_2;
wire na4455_2;
wire na4456_2;
wire na4457_2;
wire na4458_2;
wire na4459_2;
wire na4460_2;
wire na4461_2;
wire na4462_2;
wire na4463_2;
wire na4464_2;
wire na4465_2;
wire na4466_2;
wire na4467_2;
wire na4468_2;
wire na4469_2;
wire na4470_2;
wire na4471_2;
wire na4472_2;
wire na4473_2;
wire na4474_2;
wire na4475_2;
wire na4476_2;
wire na4477_2;
wire na4478_2;
wire na4479_2;
wire na4480_2;
wire na4481_2;
wire na4482_2;
wire na4483_2;
wire na4484_2;
wire na4485_2;
wire na4486_2;
wire na4487_2;
wire na4488_2;
wire na4489_2;
wire na4490_2;
wire na4491_2;
wire na4492_2;
wire na4493_2;
wire na4494_2;
wire na4495_2;
wire na4496_2;
wire na4497_2;
wire na4498_2;
wire na4499_2;
wire na4500_2;
wire na4501_2;
wire na4502_2;
wire na4503_2;
wire na4504_2;
wire na4505_2;
wire na4506_2;
wire na4507_2;
wire na4508_2;
wire na4509_2;
wire na4510_2;
wire na4511_2;
wire na4512_2;
wire na4513_2;
wire na4514_2;
wire na4515_2;
wire na4516_2;
wire na4517_2;
wire na4518_2;
wire na4519_2;
wire na4520_2;
wire na4521_2;
wire na4522_2;
wire na4523_2;
wire na4524_2;
wire na4525_2;
wire na4526_2;
wire na4527_2;
wire na4528_2;
wire na4529_2;
wire na4530_2;
wire na4531_2;
wire na4532_2;
wire na4533_2;
wire na4534_2;
wire na4535_2;
wire na4536_2;
wire na4537_2;
wire na4538_2;
wire na4539_2;
wire na4540_2;
wire na4541_2;
wire na4542_2;
wire na4543_2;
wire na4544_2;
wire na4545_2;
wire na4546_2;
wire na4547_2;
wire na4548_2;
wire na4549_2;
wire na4550_2;
wire na4551_2;
wire na4552_2;
wire na4553_2;
wire na4554_2;
wire na4555_2;
wire na4556_2;
wire na4557_2;
wire na4558_2;
wire na4559_2;
wire na4560_2;
wire na4561_2;
wire na4562_2;
wire na4563_2;
wire na4564_2;
wire na4565_2;
wire na4566_2;
wire na4567_2;
wire na4568_2;
wire na4569_2;
wire na4570_2;
wire na4571_2;
wire na4572_2;
wire na4573_2;
wire na4574_2;
wire na4575_2;
wire na4576_2;
wire na4577_2;
wire na4578_2;
wire na4579_2;
wire na4580_2;
wire na4581_2;
wire na4582_2;
wire na4583_2;
wire na4584_2;
wire na4585_2;
wire na4586_2;
wire na4587_2;
wire na4588_2;
wire na4589_2;
wire na4590_2;
wire na4591_2;
wire na4592_2;
wire na4593_2;
wire na4594_2;
wire na4595_2;
wire na4596_2;
wire na4597_2;
wire na4598_2;
wire na4599_2;
wire na4600_2;
wire na4601_2;
wire na4602_2;
wire na4603_2;
wire na4604_2;
wire na4605_2;
wire na4606_2;
wire na4607_2;
wire na4608_2;
wire na4609_2;
wire na4610_2;
wire na4611_2;
wire na4612_2;
wire na4613_2;
wire na4614_2;
wire na4615_2;
wire na4616_2;
wire na4617_2;
wire na4618_2;
wire na4619_2;
wire na4620_2;
wire na4621_2;
wire na4622_2;
wire na4623_2;
wire na4624_2;
wire na4625_2;
wire na4626_2;
wire na4627_2;
wire na4628_2;
wire na4629_2;
wire na4630_2;
wire na4631_2;
wire na4632_2;
wire na3223_93;
wire na3223_94;
wire na3223_95;
wire na3223_96;
wire na3223_97;
wire na3223_98;
wire na3223_99;
wire na3224_10;
wire na3225_93;
wire na3225_94;
wire na3225_95;
wire na3225_96;
wire na3225_97;
wire na3225_98;
wire na3225_99;
wire na3226_93;
wire na3226_94;
wire na3226_95;
wire na3226_96;
wire na3226_97;
wire na3226_98;
wire na3226_99;
wire na3227_10;
wire na3232_10;
wire na3236_10;
wire na3238_10;
wire na3240_10;
wire na3244_10;
wire na3250_10;
wire na3253_10;
wire na3261_10;
wire na3265_10;
wire na3269_10;
wire na3273_10;
wire na3280_10;
wire na3286_10;
wire na3291_10;
wire na3294_10;
wire na3297_10;
wire na3300_10;
wire na3306_10;
wire na3309_10;
wire na3314_10;
wire na3318_10;
wire na3320_10;
wire na3323_10;
wire na3326_10;
wire na3332_10;
wire na3337_10;
wire na3340_10;
wire na3345_10;
wire na3349_10;
wire na3351_10;
wire na3353_10;
wire na3355_10;
wire na3357_10;
wire na3359_10;
wire na3361_10;
wire na3363_10;
wire na3365_10;
wire na3367_10;
wire na3369_10;
wire na3371_10;
wire na3373_10;
wire na3375_10;
wire na3377_10;
wire na3379_10;
wire na3381_10;
wire na3383_10;
wire na3385_10;
wire na3387_10;
wire na3389_10;
wire na3391_10;
wire na3393_10;
wire na3395_10;
wire na3397_10;
wire na3399_10;
wire na3401_10;
wire na3403_10;
wire na3405_10;
wire na3407_10;
wire na3409_10;
wire na3411_10;
wire na3446_10;
wire na3449_10;
wire na3454_10;
wire na3456_10;
wire na3468_10;
wire na3473_10;
wire na3475_10;
wire na3477_10;
wire na3479_10;
wire na3481_10;
wire na3483_10;
wire na3485_10;
wire na3487_10;
wire na3489_10;
wire na3491_10;
wire na3493_10;
wire na3495_10;
wire na3497_10;
wire na3499_10;
wire na3501_10;
wire na3503_10;
wire na3505_10;
wire na3507_10;
wire na3509_10;
wire na3511_10;
wire na3513_10;
wire na3515_10;
wire na3517_10;
wire na3519_10;
wire na3521_10;
wire na3523_10;
wire na3533_10;
wire na3534_10;
wire na3535_10;
wire na3537_10;
wire na3540_10;
wire na3544_10;
wire na3547_10;
wire na3550_10;
wire na3553_10;
wire na3563_10;
wire na3567_10;
wire na3569_10;
wire na3573_10;
wire na3577_10;
wire na3581_10;
wire na3584_10;
wire na3587_10;
wire na3592_10;
wire na3594_10;
wire na3596_10;
wire na3598_10;
wire na3600_10;
wire na3602_10;
wire na3604_10;
wire na3606_10;
wire na3608_10;
wire na3610_10;
wire na3612_10;
wire na3614_10;
wire na3616_10;
wire na3618_10;
wire na3620_10;
wire na3622_10;
wire na3624_10;
wire na3626_10;
wire na3628_10;
wire na3630_10;
wire na3632_10;
wire na3634_10;
wire na3636_10;
wire na3638_10;
wire na3640_10;
wire na3642_10;
wire na3644_10;
wire na3646_10;
wire na3648_10;
wire na3650_10;
wire na3652_10;
wire na3654_10;
wire na3656_10;
wire na3659_10;
wire na3663_10;
wire na3666_10;
wire na3669_10;
wire na3672_10;
wire na3684_10;
wire na3686_10;
wire na3690_10;
wire na3692_10;
wire na3699_10;
wire na3704_10;
wire na3709_10;
wire na4065_10;
wire o_uart_tx;
wire na3223_100;
wire na3223_113;
wire na3223_114;
wire na3223_115;
wire na3223_116;
wire na3223_117;
wire na3223_118;
wire na3223_119;
wire na3223_120;
wire na3225_100;
wire na3226_100;
wire na3226_113;
wire na3226_114;
wire na3226_115;
wire na3226_116;
wire na3226_117;
wire na3226_118;
wire na3226_119;
wire na3226_120;

// C_AND///AND/      x17y72     80'h00_0078_00_0000_0C88_111F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2_1 ( .OUT(na2_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na7_2), .IN6(~na3_1), .IN7(~na11_1), .IN8(~na15_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2_4 ( .OUT(na2_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na233_2), .IN4(~na420_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y68     80'h00_0018_00_0000_0C88_38FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3_1 ( .OUT(na3_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na136_1), .IN6(na4_1), .IN7(1'b1), .IN8(~na645_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x49y64     80'h00_0018_00_0000_0888_2114
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4_1 ( .OUT(na4_1), .IN1(~na2229_1), .IN2(na2228_1), .IN3(~na80_1), .IN4(~na4432_2), .IN5(~na3228_1), .IN6(~na2228_2),
                   .IN7(na332_1), .IN8(~na4511_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x33y69     80'h00_0060_00_0000_0C08_FFA4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7_4 ( .OUT(na7_2), .IN1(~na1290_1), .IN2(na237_1), .IN3(na8_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y79     80'h00_0018_00_0000_0888_1AA5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1), .IN1(~na456_1), .IN2(1'b1), .IN3(na9_1), .IN4(1'b1), .IN5(na2963_2), .IN6(1'b1), .IN7(~na9_2), .IN8(~na392_1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x50y83     80'h00_0078_00_0000_0C88_411F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a9_1 ( .OUT(na9_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2962_1), .IN6(~na2965_2), .IN7(~na4570_2),
                   .IN8(na518_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a9_4 ( .OUT(na9_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na1198_1), .IN4(~na3014_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x24y71     80'h00_0018_00_0000_0C88_A4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a11_1 ( .OUT(na11_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na984_1), .IN6(na12_1), .IN7(na328_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x39y80     80'h00_0018_00_0000_0888_2141
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1), .IN1(~na1354_1), .IN2(~na232_1), .IN3(~na2713_1), .IN4(na4549_2), .IN5(~na2712_2), .IN6(~na4553_2),
                    .IN7(na1340_1), .IN8(~na3230_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x30y70     80'h00_0060_00_0000_0C08_FFC2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a15_4 ( .OUT(na15_2), .IN1(na157_1), .IN2(~na690_1), .IN3(1'b1), .IN4(na16_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x32y64     80'h00_0018_00_0000_0888_5A25
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a16_1 ( .OUT(na16_1), .IN1(~na266_1), .IN2(1'b1), .IN3(na17_1), .IN4(~na4442_2), .IN5(na2479_2), .IN6(1'b1), .IN7(~na17_2),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x28y61     80'h00_0078_00_0000_0C88_4155
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a17_1 ( .OUT(na17_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4528_2), .IN6(~na2478_1), .IN7(~na2481_2),
                    .IN8(na124_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a17_4 ( .OUT(na17_2), .IN1(~na886_1), .IN2(1'b1), .IN3(~na2529_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y71     80'h00_0018_00_0000_0C88_C2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a19_1 ( .OUT(na19_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na21_1), .IN6(~na508_2), .IN7(1'b1), .IN8(na396_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x57y69     80'h00_0018_00_0000_0888_F423
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a21_1 ( .OUT(na21_1), .IN1(1'b1), .IN2(~na22_2), .IN3(na1991_1), .IN4(~na1443_2), .IN5(~na987_1), .IN6(na22_1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x61y72     80'h00_0078_00_0000_0C88_4155
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4489_2), .IN6(~na1993_2), .IN7(~na4488_2),
                    .IN8(na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a22_4 ( .OUT(na22_2), .IN1(~na525_1), .IN2(1'b1), .IN3(~na2041_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x15y68     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a24_1 ( .OUT(na24_1), .IN1(1'b1), .IN2(na4143_2), .IN3(1'b0), .IN4(1'b0), .IN5(na4473_2), .IN6(na1617_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x25y72     80'h00_0060_00_0000_0C08_FFEC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a25_4 ( .OUT(na25_2), .IN1(1'b0), .IN2(na2_1), .IN3(na19_1), .IN4(na26_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x20y70     80'h00_0018_00_0000_0C88_C1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a26_1 ( .OUT(na26_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na28_1), .IN6(~na4071_2), .IN7(1'b1), .IN8(na27_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x26y68     80'h00_0078_00_0000_0C88_3C55
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4_1), .IN7(1'b1), .IN8(~na645_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a27_4 ( .OUT(na27_2), .IN1(~na408_1), .IN2(1'b1), .IN3(~na407_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x25y65     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a28_1 ( .OUT(na28_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na690_1), .IN7(1'b1), .IN8(na16_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x37y80     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a30_1 ( .OUT(na30_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na4074_2), .IN6(na59_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a30_2 ( .OUT(na30_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na30_1_i) );
// C_///AND/      x49y83     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a31_4 ( .OUT(na31_2), .IN1(1'b1), .IN2(na4424_2), .IN3(~na115_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x23y74     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a32_1 ( .OUT(na32_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na242_1), .IN6(na32_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a32_2 ( .OUT(na32_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na32_1_i) );
// C_AND////      x33y70     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a33_1 ( .OUT(na33_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na333_1), .IN6(1'b1), .IN7(1'b1), .IN8(na4432_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x39y74     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a34_1 ( .OUT(na34_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na39_1), .IN6(na34_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a34_2 ( .OUT(na34_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na34_1_i) );
// C_MX4b/D///      x25y76     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a35_1 ( .OUT(na35_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na53_1), .IN6(na35_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a35_2 ( .OUT(na35_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na35_1_i) );
// C_MX4b/D///      x29y67     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na36_1), .IN6(na37_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a36_2 ( .OUT(na36_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na36_1_i) );
// C_MX4b/D///      x29y72     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a37_1 ( .OUT(na37_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na51_1), .IN6(na37_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a37_2 ( .OUT(na37_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na37_1_i) );
// C_AND/D//AND/D      x66y77     80'h00_FE00_80_0000_0C88_4F88
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a38_1 ( .OUT(na38_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1149_2), .IN8(na1645_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a38_2 ( .OUT(na38_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na38_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a38_4 ( .OUT(na38_2_i), .IN1(na360_1), .IN2(na58_1), .IN3(na38_1), .IN4(na4180_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a38_5 ( .OUT(na38_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na38_2_i) );
// C_MX4b/D///      x37y73     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_1 ( .OUT(na39_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na39_1), .IN6(na40_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a39_2 ( .OUT(na39_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na39_1_i) );
// C_MX4b/D///      x35y76     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a40_1 ( .OUT(na40_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na4079_2), .IN6(na41_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a40_2 ( .OUT(na40_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na40_1_i) );
// C_MX4b/D///      x35y74     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a41_1 ( .OUT(na41_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na42_1), .IN6(na41_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a41_2 ( .OUT(na41_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na41_1_i) );
// C_MX4b/D///      x37y75     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a42_1 ( .OUT(na42_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na42_1), .IN6(na43_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a42_2 ( .OUT(na42_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na42_1_i) );
// C_MX4b/D///      x33y78     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a43_1 ( .OUT(na43_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1187_1), .IN6(na43_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a43_2 ( .OUT(na43_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na43_1_i) );
// C_MX4b/D///      x45y78     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a44_1 ( .OUT(na44_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na45_1), .IN6(na44_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a44_2 ( .OUT(na44_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na44_1_i) );
// C_MX4b/D///      x43y75     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na45_1), .IN6(na34_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a45_2 ( .OUT(na45_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na45_1_i) );
// C_MX4b/D///      x56y86     80'h00_FE00_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a46_1 ( .OUT(na46_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4081_2),
                    .IN8(na46_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a46_2 ( .OUT(na46_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na46_1_i) );
// C_MX4b/D///      x45y86     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a47_1 ( .OUT(na47_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na48_1), .IN6(na47_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a47_2 ( .OUT(na47_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na47_1_i) );
// C_MX4b/D///      x47y79     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a48_1 ( .OUT(na48_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na48_1), .IN6(na49_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a48_2 ( .OUT(na48_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na48_1_i) );
// C_MX4b/D///      x47y78     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a49_1 ( .OUT(na49_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1339_1), .IN6(na49_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a49_2 ( .OUT(na49_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na49_1_i) );
// C_MX4b/D///      x64y78     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a50_1 ( .OUT(na50_1_i), .IN1(1'b1), .IN2(~na4424_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na115_1),
                    .IN8(na50_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a50_2 ( .OUT(na50_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na50_1_i) );
// C_MX4b/D///      x23y75     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a51_1 ( .OUT(na51_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4082_2), .IN8(na52_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a51_2 ( .OUT(na51_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na51_1_i) );
// C_MX4b/D///      x26y78     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a52_1 ( .OUT(na52_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na311_1), .IN8(na52_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a52_2 ( .OUT(na52_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na52_1_i) );
// C_MX4b/D///      x21y75     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a53_1 ( .OUT(na53_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4083_2), .IN8(na112_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a53_2 ( .OUT(na53_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na53_1_i) );
// C_///AND/      x62y54     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a54_4 ( .OUT(na54_2), .IN1(1'b1), .IN2(na1451_1), .IN3(1'b1), .IN4(na55_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x56y64     80'h00_0078_00_0000_0C88_C51F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na31_2), .IN6(1'b1), .IN7(1'b1), .IN8(na56_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a55_4 ( .OUT(na55_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na528_1), .IN4(~na55_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x58y74     80'h00_FE00_00_0000_0788_5FB5
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a56_1 ( .OUT(na56_1_i), .IN1(~na31_2), .IN2(1'b0), .IN3(na4428_2), .IN4(~na56_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1149_2),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a56_2 ( .OUT(na56_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na56_1_i) );
// C_MX4b/D///      x59y80     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a57_1 ( .OUT(na57_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na4085_2), .IN6(na103_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a57_2 ( .OUT(na57_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na57_1_i) );
// C_MX4b/D///      x59y82     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a58_1 ( .OUT(na58_1_i), .IN1(1'b1), .IN2(~na4424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na4085_2), .IN6(na58_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a58_2 ( .OUT(na58_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na58_1_i) );
// C_MX4b/D///      x35y80     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a59_1 ( .OUT(na59_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na60_1), .IN6(na59_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a59_2 ( .OUT(na59_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na59_1_i) );
// C_MX4b/D///      x31y77     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a60_1 ( .OUT(na60_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na60_1), .IN6(na61_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a60_2 ( .OUT(na60_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na60_1_i) );
// C_MX4b/D///      x31y78     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a61_1 ( .OUT(na61_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na62_1), .IN6(na61_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a61_2 ( .OUT(na61_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na61_1_i) );
// C_MX4b/D///      x33y79     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a62_1 ( .OUT(na62_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na62_1), .IN6(na63_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a62_2 ( .OUT(na62_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na62_1_i) );
// C_MX4b/D///      x33y80     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a63_1 ( .OUT(na63_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na64_1), .IN6(na63_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a63_2 ( .OUT(na63_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na63_1_i) );
// C_MX4b/D///      x35y79     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a64_1 ( .OUT(na64_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na64_1), .IN6(na65_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a64_2 ( .OUT(na64_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na64_1_i) );
// C_MX4b/D///      x35y78     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a65_1 ( .OUT(na65_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1036_1), .IN6(na65_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a65_2 ( .OUT(na65_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na65_1_i) );
// C_MX4b/D///      x31y76     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a66_1 ( .OUT(na66_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na4087_2), .IN6(na66_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a66_2 ( .OUT(na66_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na66_1_i) );
// C_MX4b/D///      x31y74     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_1 ( .OUT(na67_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na68_1), .IN6(na67_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a67_2 ( .OUT(na67_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na67_1_i) );
// C_MX4b/D///      x33y73     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a68_1 ( .OUT(na68_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na68_1), .IN6(na69_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a68_2 ( .OUT(na68_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na68_1_i) );
// C_MX4b/D///      x33y74     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a69_1 ( .OUT(na69_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na4088_2), .IN6(na69_1), .IN7(1'b0),
                    .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a69_2 ( .OUT(na69_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na69_1_i) );
// C_MX4b/D///      x36y77     80'h00_FE00_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a70_1 ( .OUT(na70_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na70_1), .IN8(na71_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a70_2 ( .OUT(na70_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na70_1_i) );
// C_MX4b/D///      x36y80     80'h00_FE00_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a71_1 ( .OUT(na71_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na72_1), .IN8(na71_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a71_2 ( .OUT(na71_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na71_1_i) );
// C_MX4b/D///      x38y79     80'h00_FE00_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a72_1 ( .OUT(na72_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na72_1), .IN8(na73_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a72_2 ( .OUT(na72_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na72_1_i) );
// C_MX4b/D///      x40y82     80'h00_FE00_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a73_1 ( .OUT(na73_1_i), .IN1(~na31_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na811_1), .IN8(na73_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a73_2 ( .OUT(na73_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na73_1_i) );
// C_AND/D///      x69y88     80'h00_FE00_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1694_1), .IN6(1'b1), .IN7(~na115_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a75_2 ( .OUT(na75_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na75_1_i) );
// C_AND/D//AND/D      x68y88     80'h00_FE00_80_0000_0C88_5A1F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a76_1 ( .OUT(na76_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1694_2), .IN6(1'b1), .IN7(~na115_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a76_2 ( .OUT(na76_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na76_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a76_4 ( .OUT(na76_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na115_1), .IN4(~na76_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a76_5 ( .OUT(na76_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na76_2_i) );
// C_AND/D//AND/D      x68y84     80'h00_FE00_80_0000_0C88_5C5C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1696_2), .IN7(~na115_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a78_2 ( .OUT(na78_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a78_4 ( .OUT(na78_2_i), .IN1(1'b1), .IN2(na1696_1), .IN3(~na115_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a78_5 ( .OUT(na78_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_2_i) );
// C_AND/D//ORAND*/D      x68y82     80'h00_FE00_80_0000_0C87_5A3D
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a79_1 ( .OUT(na79_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1698_1), .IN6(1'b1), .IN7(~na115_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a79_2 ( .OUT(na79_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na79_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a79_4 ( .OUT(na79_2_i), .IN1(~na1445_2), .IN2(na1986_2), .IN3(1'b0), .IN4(~na79_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a79_5 ( .OUT(na79_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na79_2_i) );
// C_AND/D///      x58y65     80'h00_FE00_00_0000_0888_241C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1_i), .IN1(1'b1), .IN2(na81_1), .IN3(~na80_1), .IN4(~na4366_2), .IN5(~na3228_1), .IN6(na285_2), .IN7(na83_2),
                    .IN8(~na4153_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a80_2 ( .OUT(na80_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na80_1_i) );
// C_AND////      x53y62     80'h00_0018_00_0000_0888_F521
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a81_1 ( .OUT(na81_1), .IN1(~na2229_1), .IN2(~na2228_2), .IN3(na332_1), .IN4(~na4432_2), .IN5(~na2229_2), .IN6(1'b1), .IN7(1'b1),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x52y75     80'h00_0060_00_0000_0C08_FF8A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a83_4 ( .OUT(na83_2), .IN1(na1314_2), .IN2(1'b1), .IN3(na506_2), .IN4(na1296_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x47y44     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a84_4 ( .OUT(na84_2_i), .IN1(1'b1), .IN2(na536_2), .IN3(1'b1), .IN4(na3711_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a84_5 ( .OUT(na84_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na84_2_i) );
// C_AND/D//AND/D      x54y71     80'h00_FE00_80_0000_0C88_4F4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a85_1 ( .OUT(na85_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1149_2), .IN8(na4089_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a85_2 ( .OUT(na85_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na85_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a85_4 ( .OUT(na85_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1149_2), .IN4(na54_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a85_5 ( .OUT(na85_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na85_2_i) );
// C_AND/D///      x68y47     80'h00_FE00_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a87_1 ( .OUT(na87_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1639_1), .IN7(1'b1), .IN8(~na54_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a87_2 ( .OUT(na87_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na87_1_i) );
// C_AND/D//AND/D      x65y50     80'h00_FE00_80_0000_0C88_3C33
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a88_1 ( .OUT(na88_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1639_2), .IN7(1'b1), .IN8(~na54_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a88_2 ( .OUT(na88_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na88_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a88_4 ( .OUT(na88_2_i), .IN1(1'b1), .IN2(~na88_2), .IN3(1'b1), .IN4(~na54_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a88_5 ( .OUT(na88_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na88_2_i) );
// C_AND/D//AND/D      x67y52     80'h00_FE00_80_0000_0C88_3A3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1641_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na54_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a89_2 ( .OUT(na89_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a89_4 ( .OUT(na89_2_i), .IN1(na1641_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na54_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a89_5 ( .OUT(na89_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_2_i) );
// C_ORAND*////D      x61y73     80'h00_FE18_00_0000_0788_DA5D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a90_1 ( .OUT(na90_1), .IN1(~na4253_2), .IN2(na91_1), .IN3(~na85_1), .IN4(1'b0), .IN5(na4043_1), .IN6(1'b0), .IN7(~na4365_2),
                    .IN8(na98_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a90_5 ( .OUT(na90_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na90_1) );
// C_ORAND////      x69y52     80'h00_0018_00_0000_0C88_3DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a91_1 ( .OUT(na91_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na987_1), .IN6(na4092_2), .IN7(1'b0), .IN8(~na92_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x70y50     80'h00_0018_00_0000_0C88_2CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a92_1 ( .OUT(na92_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1451_1), .IN7(na93_1), .IN8(~na55_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x68y61     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_1 ( .OUT(na93_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na525_1), .IN6(1'b1), .IN7(~na2041_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x65y76     80'h00_0078_00_0000_0C88_AA3A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a94_1 ( .OUT(na94_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na95_1), .IN6(1'b1), .IN7(na598_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a94_4 ( .OUT(na94_2), .IN1(na534_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na78_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x67y73     80'h00_0078_00_0000_0C88_C1C8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a95_1 ( .OUT(na95_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4489_2), .IN6(~na1993_2), .IN7(1'b1), .IN8(na1990_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a95_4 ( .OUT(na95_2), .IN1(na4489_2), .IN2(na1993_2), .IN3(1'b1), .IN4(na612_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x66y74     80'h00_0018_00_0040_0A2B_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a98_1 ( .OUT(na98_1), .IN1(1'b1), .IN2(~na1993_2), .IN3(1'b1), .IN4(~na1990_1), .IN5(1'b1), .IN6(~na3241_2), .IN7(1'b0),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x61y78     80'h00_FE00_00_0040_0A3C_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_1 ( .OUT(na103_1_i), .IN1(1'b1), .IN2(~na4424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na4148_2), .IN6(na103_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a103_2 ( .OUT(na103_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na103_1_i) );
// C_MX4b/D///      x62y74     80'h00_FE00_00_0040_0AC8_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a104_1 ( .OUT(na104_1_i), .IN1(na105_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4094_2),
                     .IN8(~na104_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a104_2 ( .OUT(na104_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na104_1_i) );
// C_ORAND/D///      x63y75     80'h00_FE00_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a105_1 ( .OUT(na105_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na105_1), .IN6(na4090_2), .IN7(1'b0), .IN8(na3243_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a105_2 ( .OUT(na105_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na105_1_i) );
// C_MX4b/D///      x58y75     80'h00_FE00_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a107_1 ( .OUT(na107_1_i), .IN1(na105_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na107_1),
                     .IN8(na1628_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a107_2 ( .OUT(na107_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na107_1_i) );
// C_MX4b/D///      x62y76     80'h00_FE00_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a108_1 ( .OUT(na108_1_i), .IN1(~na105_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1630_2),
                     .IN8(na108_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a108_2 ( .OUT(na108_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na108_1_i) );
// C_MX4b/D///      x59y75     80'h00_FE00_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a109_1 ( .OUT(na109_1_i), .IN1(na105_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4097_2),
                     .IN8(na1628_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a109_2 ( .OUT(na109_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na109_1_i) );
// C_MX4b/D///      x20y64     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a110_1 ( .OUT(na110_1_i), .IN1(1'b1), .IN2(~na1487_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1369_1),
                     .IN8(na110_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a110_2 ( .OUT(na110_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na110_1_i) );
// C_MX4b/D///      x23y76     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a111_1 ( .OUT(na111_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na118_1), .IN6(na111_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a111_2 ( .OUT(na111_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na111_1_i) );
// C_MX4b/D///      x28y74     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a112_1 ( .OUT(na112_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na4099_2), .IN6(na111_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a112_2 ( .OUT(na112_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na112_1_i) );
// C_MX4b/D///      x15y66     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a113_1 ( .OUT(na113_1_i), .IN1(1'b1), .IN2(~na1487_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na4098_2), .IN6(na113_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a113_2 ( .OUT(na113_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na113_1_i) );
// C_MX4b/D///      x21y63     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a114_1 ( .OUT(na114_1_i), .IN1(1'b1), .IN2(na1487_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na114_1), .IN6(na113_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a114_2 ( .OUT(na114_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na114_1_i) );
// C_MX4b/D///      x68y79     80'h00_FE00_00_0040_0A51_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a115_1 ( .OUT(na115_1_i), .IN1(na4078_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4103_2), .IN5(~na117_1), .IN6(1'b0), .IN7(na115_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a115_2 ( .OUT(na115_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na115_1_i) );
// C_AND///AND/      x69y75     80'h00_0078_00_0000_0C88_433A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a117_1 ( .OUT(na117_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na94_1), .IN7(~na603_2), .IN8(na98_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a117_4 ( .OUT(na117_2), .IN1(na90_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na50_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x25y75     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a118_1 ( .OUT(na118_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na118_1), .IN6(na127_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a118_2 ( .OUT(na118_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na118_1_i) );
// C_MX4b/D///      x15y76     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a119_1 ( .OUT(na119_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na125_1), .IN6(na119_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a119_2 ( .OUT(na119_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na119_1_i) );
// C_///AND/      x15y74     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a120_4 ( .OUT(na120_2), .IN1(1'b1), .IN2(~na299_1), .IN3(1'b1), .IN4(na4442_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x25y53     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a121_4 ( .OUT(na121_2), .IN1(1'b1), .IN2(na122_1), .IN3(1'b1), .IN4(na1495_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x19y48     80'h00_0078_00_0000_0C88_A3F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a122_1 ( .OUT(na122_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na120_2), .IN7(na123_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a122_4 ( .OUT(na122_2), .IN1(~na196_2), .IN2(~na122_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*/D///      x18y63     80'h00_FE00_00_0000_0788_5FD3
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a123_1 ( .OUT(na123_1_i), .IN1(1'b0), .IN2(~na120_2), .IN3(~na123_1), .IN4(na1495_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na1149_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a123_2 ( .OUT(na123_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na123_1_i) );
// C_MX4b/D///      x20y60     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a124_1 ( .OUT(na124_1_i), .IN1(1'b1), .IN2(na1487_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na4105_2), .IN6(na299_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a124_2 ( .OUT(na124_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na124_1_i) );
// C_MX4b/D///      x13y77     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a125_1 ( .OUT(na125_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na125_1), .IN6(na126_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a125_2 ( .OUT(na125_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na125_1_i) );
// C_MX4b/D///      x17y70     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a126_1 ( .OUT(na126_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na1367_1), .IN6(na126_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a126_2 ( .OUT(na126_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na126_1_i) );
// C_MX4b/D///      x25y74     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a127_1 ( .OUT(na127_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na128_1), .IN6(na127_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a127_2 ( .OUT(na127_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na127_1_i) );
// C_MX4b/D///      x25y73     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na128_1), .IN6(na4106_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a128_2 ( .OUT(na128_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na128_1_i) );
// C_MX4b/D///      x27y71     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a129_1 ( .OUT(na129_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na129_1), .IN6(na32_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a129_2 ( .OUT(na129_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na129_1_i) );
// C_MX4b/D///      x17y66     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a130_1 ( .OUT(na130_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na131_1), .IN6(na130_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a130_2 ( .OUT(na130_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na130_1_i) );
// C_MX4b/D///      x17y67     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a131_1 ( .OUT(na131_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na131_1), .IN6(na132_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a131_2 ( .OUT(na131_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na131_1_i) );
// C_MX4b/D///      x19y70     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a132_1 ( .OUT(na132_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na133_1), .IN6(na132_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a132_2 ( .OUT(na132_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na132_1_i) );
// C_MX4b/D///      x17y75     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a133_1 ( .OUT(na133_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4107_2),
                     .IN8(na1365_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a133_2 ( .OUT(na133_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na133_1_i) );
// C_MX4b/D///      x18y83     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a134_1 ( .OUT(na134_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na134_1),
                     .IN8(na135_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a134_2 ( .OUT(na134_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na134_1_i) );
// C_MX4b/D///      x18y84     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a135_1 ( .OUT(na135_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na153_1), .IN6(na4108_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a135_2 ( .OUT(na135_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na135_1_i) );
// C_MX4b/D///      x21y69     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a136_1 ( .OUT(na136_1_i), .IN1(1'b1), .IN2(na137_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na136_1), .IN6(na3147_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a136_2 ( .OUT(na136_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na136_1_i) );
// C_///AND/      x33y70     80'h00_0060_00_0000_0C08_FF53
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a137_4 ( .OUT(na137_2), .IN1(1'b1), .IN2(~na138_1), .IN3(~na139_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x27y68     80'h00_0018_00_0000_0888_CD35
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(~na28_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na27_1), .IN5(~na21_1), .IN6(na508_2), .IN7(1'b0), .IN8(na27_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y75     80'h00_0018_00_0000_0888_3582
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a139_1 ( .OUT(na139_1), .IN1(na3246_1), .IN2(~na146_1), .IN3(na506_2), .IN4(na3248_1), .IN5(~na143_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(~na3249_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x41y69     80'h00_0018_00_0000_0888_4CC8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a143_1 ( .OUT(na143_1), .IN1(na145_1), .IN2(na690_1), .IN3(1'b1), .IN4(na4154_2), .IN5(1'b1), .IN6(na900_1), .IN7(~na4152_2),
                     .IN8(na16_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x47y75     80'h00_0018_00_0000_0C88_85FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a145_1 ( .OUT(na145_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1314_2), .IN6(1'b1), .IN7(na506_2), .IN8(na1296_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x53y70     80'h00_0018_00_0000_0888_28F8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a146_1 ( .OUT(na146_1), .IN1(na145_1), .IN2(na508_2), .IN3(1'b1), .IN4(1'b1), .IN5(na21_1), .IN6(na285_1), .IN7(na551_1),
                     .IN8(~na4154_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x19y83     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a153_1 ( .OUT(na153_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na153_1), .IN6(na154_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a153_2 ( .OUT(na153_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na153_1_i) );
// C_MX4b/D///      x19y84     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a154_1 ( .OUT(na154_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na1364_1), .IN6(na154_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a154_2 ( .OUT(na154_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na154_1_i) );
// C_///ORAND/      x13y64     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a155_4 ( .OUT(na155_2), .IN1(~na1614_1), .IN2(~na405_2), .IN3(~na4474_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x14y68     80'h00_0018_00_0000_0C88_37FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a156_1 ( .OUT(na156_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4470_2), .IN6(~na2_2), .IN7(1'b0), .IN8(~na1610_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x19y73     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a157_1 ( .OUT(na157_1_i), .IN1(1'b1), .IN2(na137_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na157_1), .IN6(na3148_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a157_2 ( .OUT(na157_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na157_1_i) );
// C_MX4b/D///      x19y86     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a158_1 ( .OUT(na158_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4112_2),
                     .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a158_2 ( .OUT(na158_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na158_1_i) );
// C_MX4b/D///      x20y84     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a159_1 ( .OUT(na159_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4113_2),
                     .IN8(na159_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a159_2 ( .OUT(na159_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na159_1_i) );
// C_MX4b/D///      x17y83     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a160_1 ( .OUT(na160_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na160_1), .IN6(na161_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a160_2 ( .OUT(na160_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na160_1_i) );
// C_MX4b/D///      x19y82     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a161_1 ( .OUT(na161_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na1357_1), .IN6(na161_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a161_2 ( .OUT(na161_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na161_1_i) );
// C_MX4b/D///      x38y68     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a162_1 ( .OUT(na162_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4170_2),
                     .IN8(na162_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a162_2 ( .OUT(na162_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na162_1_i) );
// C_MX4b/D///      x13y83     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a163_1 ( .OUT(na163_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na164_1), .IN6(na4114_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a163_2 ( .OUT(na163_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na163_1_i) );
// C_MX4b/D///      x17y81     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a164_1 ( .OUT(na164_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na164_1), .IN6(na4115_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a164_2 ( .OUT(na164_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na164_1_i) );
// C_MX4b/D///      x17y82     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a165_1 ( .OUT(na165_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na167_1), .IN6(na165_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a165_2 ( .OUT(na165_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na165_1_i) );
// C_MX4b/D///      x17y79     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a166_1 ( .OUT(na166_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na166_1), .IN6(na165_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a166_2 ( .OUT(na166_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na166_1_i) );
// C_MX4b/D///      x15y77     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a167_1 ( .OUT(na167_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na1355_1), .IN6(na4116_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a167_2 ( .OUT(na167_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na167_1_i) );
// C_MX4b/D///      x15y80     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a168_1 ( .OUT(na168_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na4118_2), .IN6(na168_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a168_2 ( .OUT(na168_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na168_1_i) );
// C_MX4b/D///      x17y77     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a169_1 ( .OUT(na169_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na169_1), .IN6(na168_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a169_2 ( .OUT(na169_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na169_1_i) );
// C_MX4b/D///      x16y80     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a170_1 ( .OUT(na170_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na171_1),
                     .IN8(na170_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a170_2 ( .OUT(na170_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na170_1_i) );
// C_MX4b/D///      x16y77     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a171_1 ( .OUT(na171_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na171_1),
                     .IN8(na174_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a171_2 ( .OUT(na171_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na171_1_i) );
// C_AND/D///      x13y47     80'h00_FE00_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a173_1 ( .OUT(na173_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na299_1), .IN7(na1688_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a173_2 ( .OUT(na173_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na173_1_i) );
// C_MX4b/D///      x16y76     80'h00_FE00_00_0040_0AC4_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a174_1 ( .OUT(na174_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na175_1),
                     .IN8(na174_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a174_2 ( .OUT(na174_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na174_1_i) );
// C_MX2a////      x16y71     80'h00_0018_00_0040_0CCC_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a175_1 ( .OUT(na175_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na176_2), .IN4(~na187_2), .IN5(~na1370_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x20y69     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a176_4 ( .OUT(na176_2), .IN1(1'b1), .IN2(1'b1), .IN3(na123_1), .IN4(na3252_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x14y64     80'h00_0018_00_0000_0C88_DCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a178_1 ( .OUT(na178_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na119_1), .IN7(~na179_1), .IN8(na3254_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x18y59     80'h00_0018_00_0040_0C92_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a179_1 ( .OUT(na179_1), .IN1(1'b1), .IN2(na2478_1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b1), .IN6(~na2478_2), .IN7(1'b1), .IN8(na4525_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x15y64     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a180_1 ( .OUT(na180_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3255_1), .IN6(1'b0), .IN7(na4582_2), .IN8(~na2499_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x17y57     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a181_1 ( .OUT(na181_1), .IN1(na182_1), .IN2(1'b1), .IN3(1'b1), .IN4(na214_2), .IN5(na832_1), .IN6(na827_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x21y55     80'h00_0018_00_0000_0C88_12FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_1 ( .OUT(na182_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2479_2), .IN6(~na2477_1), .IN7(~na4529_2),
                     .IN8(~na4527_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x20y72     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a187_4 ( .OUT(na187_2), .IN1(na1484_2), .IN2(na119_1), .IN3(1'b0), .IN4(na188_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x16y66     80'h00_0018_00_0000_0C88_2CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a188_1 ( .OUT(na188_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na113_1), .IN7(na189_2), .IN8(~na214_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x16y63     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a189_4 ( .OUT(na189_2), .IN1(~na216_1), .IN2(1'b1), .IN3(~na4134_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D//AND/D      x16y50     80'h00_FE00_80_0000_0C88_A333
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a190_1 ( .OUT(na190_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na299_1), .IN7(na1688_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a190_2 ( .OUT(na190_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na190_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a190_4 ( .OUT(na190_2_i), .IN1(1'b1), .IN2(~na299_1), .IN3(1'b1), .IN4(~na190_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a190_5 ( .OUT(na190_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na190_2_i) );
// C_AND/D//AND/D      x15y51     80'h00_FE00_80_0000_0C88_C3C3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a192_1 ( .OUT(na192_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na299_1), .IN7(1'b1), .IN8(na1690_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a192_2 ( .OUT(na192_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na192_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a192_4 ( .OUT(na192_2_i), .IN1(1'b1), .IN2(~na299_1), .IN3(1'b1), .IN4(na1690_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a192_5 ( .OUT(na192_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na192_2_i) );
// C_AND/D//ORAND*/D      x15y50     80'h00_FE00_80_0000_0C87_A33D
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a193_1 ( .OUT(na193_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na299_1), .IN7(na1692_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a193_2 ( .OUT(na193_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na193_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a193_4 ( .OUT(na193_2_i), .IN1(~na4444_2), .IN2(na2474_2), .IN3(1'b0), .IN4(~na4121_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a193_5 ( .OUT(na193_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na193_2_i) );
// C_ORAND////      x25y44     80'h00_0018_00_0000_0888_FE3A
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a194_1 ( .OUT(na194_1), .IN1(na3259_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1495_2), .IN5(na196_2), .IN6(na122_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x21y59     80'h00_0060_00_0000_0C08_FF21
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a196_4 ( .OUT(na196_2), .IN1(~na886_1), .IN2(~na4542_2), .IN3(na17_1), .IN4(~na4442_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x24y50     80'h00_FE00_00_0000_0C88_38FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a197_1 ( .OUT(na197_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na210_1), .IN6(na209_1), .IN7(1'b1), .IN8(~na208_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a197_2 ( .OUT(na197_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na197_1_i) );
// C_OR////D      x25y39     80'h00_FE18_00_0000_0EEE_0C03
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a198_1 ( .OUT(na198_1), .IN1(1'b0), .IN2(~na194_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3262_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a198_5 ( .OUT(na198_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na198_1) );
// C_AND/D//AND/D      x24y66     80'h00_FE00_80_0000_0C88_4F5A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a200_1 ( .OUT(na200_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1149_2), .IN8(na200_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a200_2 ( .OUT(na200_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na200_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a200_4 ( .OUT(na200_2_i), .IN1(na121_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a200_5 ( .OUT(na200_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na200_2_i) );
// C_///AND/D      x40y47     80'h00_FE00_80_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a201_4 ( .OUT(na201_2_i), .IN1(~na121_2), .IN2(1'b1), .IN3(na1709_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a201_5 ( .OUT(na201_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na201_2_i) );
// C_AND/D///      x25y38     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a202_1 ( .OUT(na202_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4124_2), .IN7(1'b1), .IN8(na3525_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a202_2 ( .OUT(na202_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na202_1_i) );
// C_AND////D      x30y42     80'h00_FE18_00_0000_0888_53FC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a203_1 ( .OUT(na203_1), .IN1(1'b1), .IN2(na204_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na204_1), .IN7(~na201_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a203_5 ( .OUT(na203_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na203_1) );
// C_AND/D//AND/D      x39y48     80'h00_FE00_80_0000_0C88_A5F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a204_1 ( .OUT(na204_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na121_2), .IN6(1'b1), .IN7(na1709_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a204_2 ( .OUT(na204_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na204_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a204_4 ( .OUT(na204_2_i), .IN1(~na121_2), .IN2(~na204_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a204_5 ( .OUT(na204_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na204_2_i) );
// C_///AND/D      x27y46     80'h00_FE00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a205_4 ( .OUT(na205_2_i), .IN1(na4125_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3525_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a205_5 ( .OUT(na205_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na205_2_i) );
// C_AND/D//AND/D      x41y44     80'h00_FE00_80_0000_0C88_C5C5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a207_1 ( .OUT(na207_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na121_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1711_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a207_2 ( .OUT(na207_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na207_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a207_4 ( .OUT(na207_2_i), .IN1(~na121_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1711_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a207_5 ( .OUT(na207_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na207_2_i) );
// C_MX4b/D///      x18y60     80'h00_FE00_00_0040_0AC8_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a208_1 ( .OUT(na208_1_i), .IN1(na212_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4128_2),
                     .IN8(~na208_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a208_2 ( .OUT(na208_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na208_1_i) );
// C_MX4b/D///      x13y62     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a209_1 ( .OUT(na209_1_i), .IN1(na212_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na4129_2), .IN6(na1714_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a209_2 ( .OUT(na209_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na209_1_i) );
// C_MX4b/D///      x15y57     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a210_1 ( .OUT(na210_1_i), .IN1(na212_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na210_1), .IN6(na1714_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a210_2 ( .OUT(na210_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na210_1_i) );
// C_MX4b/D///      x18y55     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a211_1 ( .OUT(na211_1_i), .IN1(~na212_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1716_1), .IN6(na4130_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a211_2 ( .OUT(na211_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na211_1_i) );
// C_ORAND/D///      x13y55     80'h00_FE00_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a212_1 ( .OUT(na212_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na212_1), .IN6(na4469_2), .IN7(na3263_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a212_2 ( .OUT(na212_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na212_1_i) );
// C_AND/D//AND/D      x20y62     80'h00_FE00_80_0000_0C88_4F88
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a214_1 ( .OUT(na214_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1149_2), .IN8(na1705_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a214_2 ( .OUT(na214_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na214_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a214_4 ( .OUT(na214_2_i), .IN1(na216_1), .IN2(na113_1), .IN3(na4134_2), .IN4(na214_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a214_5 ( .OUT(na214_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na214_2_i) );
// C_AND/D//AND/D      x27y63     80'h00_FE00_80_0000_0C88_2F4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a216_1 ( .OUT(na216_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1707_1), .IN8(~na4366_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a216_2 ( .OUT(na216_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na216_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a216_4 ( .OUT(na216_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1149_2), .IN4(na1705_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a216_5 ( .OUT(na216_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na216_2_i) );
// C_AND/D//AND/D      x36y82     80'h00_FE00_80_0000_0C88_5A4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a217_1 ( .OUT(na217_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na218_1), .IN6(1'b1), .IN7(~na1149_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a217_2 ( .OUT(na217_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na217_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a217_4 ( .OUT(na217_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1149_2), .IN4(na217_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a217_5 ( .OUT(na217_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na217_2_i) );
// C_AND////      x45y79     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a218_1 ( .OUT(na218_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na219_2), .IN7(na1517_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x39y72     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a219_4 ( .OUT(na219_2), .IN1(~na220_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1337_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x25y89     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a220_1 ( .OUT(na220_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na232_1), .IN7(1'b1), .IN8(~na1347_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x57y65     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a221_1 ( .OUT(na221_1_i), .IN1(na1465_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na221_1), .IN6(na330_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a221_2 ( .OUT(na221_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na221_1_i) );
// C_ORAND*////D      x37y89     80'h00_FE18_00_0000_0788_DA3D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a222_1 ( .OUT(na222_1), .IN1(~na1118_2), .IN2(na223_2), .IN3(1'b0), .IN4(~na217_2), .IN5(na1564_1), .IN6(1'b0), .IN7(~na1346_1),
                     .IN8(na229_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a222_5 ( .OUT(na222_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na222_1) );
// C_///ORAND/      x61y76     80'h00_0060_00_0000_0C08_FF5D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a223_4 ( .OUT(na223_2), .IN1(~na1354_1), .IN2(na4581_2), .IN3(~na224_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x58y81     80'h00_0018_00_0000_0C88_21FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a224_1 ( .OUT(na224_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2769_1), .IN6(~na219_2), .IN7(na1517_2),
                     .IN8(~na1050_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x35y92     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a225_4 ( .OUT(na225_2), .IN1(1'b1), .IN2(1'b1), .IN3(na226_1), .IN4(na1113_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x40y89     80'h00_0078_00_0000_0C88_528C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a226_1 ( .OUT(na226_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2712_2), .IN6(~na4553_2), .IN7(~na2713_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a226_4 ( .OUT(na226_2), .IN1(1'b1), .IN2(na4553_2), .IN3(na2713_1), .IN4(na1127_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x34y86     80'h00_0018_00_0040_0A8E_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a229_1 ( .OUT(na229_1), .IN1(na2712_2), .IN2(1'b1), .IN3(~na2713_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(~na3270_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//AND/D      x41y80     80'h00_FE00_80_0000_0C88_5E88
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a232_1 ( .OUT(na232_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na222_1), .IN6(na232_1), .IN7(~na4141_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a232_2 ( .OUT(na232_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na232_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a232_4 ( .OUT(na232_2_i), .IN1(na434_1), .IN2(na4144_2), .IN3(na432_2), .IN4(na4200_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a232_5 ( .OUT(na232_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na232_2_i) );
// C_AND///AND/      x18y69     80'h00_0078_00_0000_0C88_515C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a233_1 ( .OUT(na233_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1614_1), .IN6(~na405_2), .IN7(~na4474_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a233_4 ( .OUT(na233_2), .IN1(1'b1), .IN2(na2_1), .IN3(~na19_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x13y63     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a234_1 ( .OUT(na234_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1614_1), .IN6(1'b1), .IN7(~na4474_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x15y65     80'h00_0060_00_0000_0C08_FF31
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a235_4 ( .OUT(na235_2), .IN1(~na4471_2), .IN2(~na2_2), .IN3(1'b1), .IN4(~na1610_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x14y65     80'h00_0018_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a236_1 ( .OUT(na236_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na4472_2), .IN8(~na1610_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x21y72     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a237_1 ( .OUT(na237_1_i), .IN1(1'b1), .IN2(~na137_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na3149_1), .IN6(na237_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a237_2 ( .OUT(na237_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na237_1_i) );
// C_MX4b/D///      x32y85     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a238_1 ( .OUT(na238_1_i), .IN1(1'b1), .IN2(na232_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na238_1),
                     .IN8(na239_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a238_2 ( .OUT(na238_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na238_1_i) );
// C_MX4b/D///      x32y86     80'h00_FE00_00_0040_0AC3_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a239_1 ( .OUT(na239_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na241_1),
                     .IN8(na239_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a239_2 ( .OUT(na239_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na239_1_i) );
// C_MX4b/D///      x32y84     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a240_1 ( .OUT(na240_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na238_1),
                     .IN8(na240_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a240_2 ( .OUT(na240_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na240_1_i) );
// C_MX4b/D///      x32y83     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a241_1 ( .OUT(na241_1_i), .IN1(1'b1), .IN2(na232_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na241_1),
                     .IN8(na240_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a241_2 ( .OUT(na241_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na241_1_i) );
// C_MX4b/D///      x23y73     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a242_1 ( .OUT(na242_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na242_1), .IN6(na4146_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a242_2 ( .OUT(na242_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na242_1_i) );
// C_MX4b/D///      x27y75     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a243_1 ( .OUT(na243_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na243_1), .IN6(na244_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a243_2 ( .OUT(na243_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na243_1_i) );
// C_MX4b/D///      x29y74     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a244_1 ( .OUT(na244_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na4147_2), .IN6(na244_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a244_2 ( .OUT(na244_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na244_1_i) );
// C_MX4b/D///      x30y74     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a245_1 ( .OUT(na245_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na247_1),
                     .IN8(na245_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a245_2 ( .OUT(na245_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na245_1_i) );
// C_MX4b/D///      x60y79     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a246_1 ( .OUT(na246_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na4148_2), .IN6(na58_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a246_2 ( .OUT(na246_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na246_1_i) );
// C_MX4b/D///      x40y73     80'h00_FE00_00_0040_0AC8_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a247_1 ( .OUT(na247_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na247_1), .IN8(~na248_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a247_2 ( .OUT(na247_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na247_1_i) );
// C_MX2b////      x58y72     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a248_1 ( .OUT(na248_1), .IN1(na349_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na260_2), .IN8(~na249_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x62y68     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a249_1 ( .OUT(na249_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na326_1), .IN8(na3272_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x60y67     80'h00_0060_00_0000_0C08_FFCD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a251_4 ( .OUT(na251_2), .IN1(~na252_1), .IN2(na3274_2), .IN3(1'b0), .IN4(na327_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x61y63     80'h00_0018_00_0040_0C92_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a252_1 ( .OUT(na252_1), .IN1(1'b1), .IN2(na2228_2), .IN3(1'b0), .IN4(1'b1), .IN5(~na2229_2), .IN6(1'b1), .IN7(na2226_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x61y67     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a253_1 ( .OUT(na253_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3278_2), .IN6(~na2248_1), .IN7(1'b0), .IN8(~na3275_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x58y59     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a254_1 ( .OUT(na254_1), .IN1(1'b1), .IN2(na255_2), .IN3(1'b1), .IN4(~na4160_2), .IN5(1'b0), .IN6(1'b0), .IN7(na653_1), .IN8(na648_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y60     80'h00_0060_00_0000_0C08_FF14
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a255_4 ( .OUT(na255_2), .IN1(~na2229_2), .IN2(na2228_1), .IN3(~na2226_2), .IN4(~na4508_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x60y71     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a260_4 ( .OUT(na260_2), .IN1(1'b0), .IN2(na261_2), .IN3(na1462_2), .IN4(na327_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y70     80'h00_0060_00_0000_0C08_FFA2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a261_4 ( .OUT(na261_2), .IN1(na221_1), .IN2(~na295_1), .IN3(na262_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x54y63     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a262_1 ( .OUT(na262_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4161_2), .IN6(1'b1), .IN7(~na297_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x32y57     80'h00_FE00_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a264_1 ( .OUT(na264_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na333_1), .IN6(1'b1), .IN7(na1722_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a264_2 ( .OUT(na264_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na264_1_i) );
// C_AND/D//AND/D      x31y60     80'h00_FE00_80_0000_0C88_A5F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a265_1 ( .OUT(na265_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na333_1), .IN6(1'b1), .IN7(na1722_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a265_2 ( .OUT(na265_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na265_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a265_4 ( .OUT(na265_2_i), .IN1(~na333_1), .IN2(~na265_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a265_5 ( .OUT(na265_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na265_2_i) );
// C_AND/D///      x39y63     80'h00_FE00_00_0000_0888_4412
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a266_1 ( .OUT(na266_1_i), .IN1(na145_1), .IN2(~na285_1), .IN3(~na1149_2), .IN4(~na4442_2), .IN5(~na266_1), .IN6(na285_2),
                     .IN7(~na17_2), .IN8(na4068_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a266_2 ( .OUT(na266_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na266_1_i) );
// C_AND/D//ORAND*/D      x45y58     80'h00_FE00_80_0000_0C87_A5B3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a268_1 ( .OUT(na268_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na333_1), .IN6(1'b1), .IN7(na1726_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a268_2 ( .OUT(na268_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na268_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a268_4 ( .OUT(na268_2_i), .IN1(1'b0), .IN2(~na268_1), .IN3(na2223_2), .IN4(~na4434_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a268_5 ( .OUT(na268_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na268_2_i) );
// C_///AND/D      x48y39     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a269_4 ( .OUT(na269_2_i), .IN1(1'b1), .IN2(na273_2), .IN3(1'b1), .IN4(na3719_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a269_5 ( .OUT(na269_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na269_2_i) );
// C_AND/D//AND/D      x32y60     80'h00_FE00_80_0000_0C88_C5C5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a270_1 ( .OUT(na270_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na333_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1724_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a270_2 ( .OUT(na270_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na270_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a270_4 ( .OUT(na270_2_i), .IN1(~na333_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1724_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a270_5 ( .OUT(na270_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na270_2_i) );
// C_AND/D///      x48y39     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a272_1 ( .OUT(na272_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na273_1), .IN7(1'b1), .IN8(na3719_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a272_2 ( .OUT(na272_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na272_1_i) );
// C_AND////D      x53y38     80'h00_FE18_00_0000_0888_3CF3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a273_1 ( .OUT(na273_1), .IN1(1'b1), .IN2(~na274_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na274_2), .IN7(1'b1), .IN8(~na277_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a273_5 ( .OUT(na273_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na273_1) );
// C_AND/D//AND/D      x65y38     80'h00_FE00_80_0000_0C88_A5F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a274_1 ( .OUT(na274_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na275_2), .IN6(1'b1), .IN7(na1733_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a274_2 ( .OUT(na274_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na274_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a274_4 ( .OUT(na274_2_i), .IN1(~na275_2), .IN2(~na274_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a274_5 ( .OUT(na274_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na274_2_i) );
// C_///AND/      x57y45     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a275_4 ( .OUT(na275_2), .IN1(na1473_2), .IN2(1'b1), .IN3(na276_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y55     80'h00_0018_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a276_1 ( .OUT(na276_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na33_1), .IN7(na326_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x62y40     80'h00_FE00_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a277_1 ( .OUT(na277_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na275_2), .IN6(1'b1), .IN7(na1733_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a277_2 ( .OUT(na277_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na277_1_i) );
// C_AND/D//AND/D      x68y35     80'h00_FE00_80_0000_0C88_C5C5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a280_1 ( .OUT(na280_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na275_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1735_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a280_2 ( .OUT(na280_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na280_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a280_4 ( .OUT(na280_2_i), .IN1(~na275_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1735_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a280_5 ( .OUT(na280_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na280_2_i) );
// C_AND/D//AND/D      x49y66     80'h00_FE00_80_0000_0C88_5C5A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a281_1 ( .OUT(na281_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na281_2), .IN7(~na1149_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a281_2 ( .OUT(na281_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na281_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a281_4 ( .OUT(na281_2_i), .IN1(na275_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a281_5 ( .OUT(na281_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na281_2_i) );
// C_MX4b/D///      x46y62     80'h00_FE00_00_0040_0AC8_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a282_1 ( .OUT(na282_1_i), .IN1(1'b1), .IN2(na1383_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4151_2),
                     .IN8(~na282_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a282_2 ( .OUT(na282_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na282_1_i) );
// C_MX4b/D///      x46y63     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a283_1 ( .OUT(na283_1_i), .IN1(1'b1), .IN2(na1383_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na283_1),
                     .IN8(na1728_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a283_2 ( .OUT(na283_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na283_1_i) );
// C_MX4b/D///      x48y62     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_1 ( .OUT(na284_1_i), .IN1(1'b1), .IN2(~na1383_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1730_2),
                     .IN8(na284_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a284_2 ( .OUT(na284_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na284_1_i) );
// C_ORAND/D//ORAND/D      x51y70     80'h00_FE00_80_0000_0C88_5B5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a285_1 ( .OUT(na285_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3290_2), .IN6(~na3279_1), .IN7(~na1149_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a285_2 ( .OUT(na285_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na285_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a285_4 ( .OUT(na285_2_i), .IN1(na3290_1), .IN2(na321_1), .IN3(~na1149_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a285_5 ( .OUT(na285_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na285_2_i) );
// C_AND/D//ORAND*/D      x20y87     80'h00_FE00_80_0000_0C87_1CD5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a287_1 ( .OUT(na287_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1620_1), .IN7(~na287_2), .IN8(~na4156_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a287_2 ( .OUT(na287_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na287_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a287_4 ( .OUT(na287_2_i), .IN1(~na3700_1), .IN2(1'b0), .IN3(~na287_2), .IN4(na1296_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a287_5 ( .OUT(na287_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na287_2_i) );
// C_AND/D//AND/D      x17y86     80'h00_FE00_80_0000_0C88_5252
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a288_1 ( .OUT(na288_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1618_1), .IN6(~na288_2), .IN7(~na287_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a288_2 ( .OUT(na288_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na288_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a288_4 ( .OUT(na288_2_i), .IN1(na1626_1), .IN2(~na288_2), .IN3(~na287_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a288_5 ( .OUT(na288_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na288_2_i) );
// C_OR/D///      x14y84     80'h00_FE00_00_0000_0CEE_EC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a289_1 ( .OUT(na289_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1620_2), .IN7(na287_2), .IN8(na4158_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a289_2 ( .OUT(na289_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na289_1_i) );
// C_AND/D//AND/D      x16y88     80'h00_FE00_80_0000_0C88_5252
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a292_1 ( .OUT(na292_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1622_2), .IN6(~na288_2), .IN7(~na287_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a292_2 ( .OUT(na292_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na292_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a292_4 ( .OUT(na292_2_i), .IN1(na1622_1), .IN2(~na288_2), .IN3(~na287_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a292_5 ( .OUT(na292_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na292_2_i) );
// C_///AND/D      x17y76     80'h00_FE00_80_0000_0C08_FF1C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a293_4 ( .OUT(na293_2_i), .IN1(1'b1), .IN2(na1624_1), .IN3(~na287_2), .IN4(~na4156_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a293_5 ( .OUT(na293_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na293_2_i) );
// C_///OR/D      x16y81     80'h00_FE00_80_0000_0C0E_FFEC
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a294_4 ( .OUT(na294_2_i), .IN1(1'b0), .IN2(na1624_2), .IN3(na287_2), .IN4(na4158_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a294_5 ( .OUT(na294_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na294_2_i) );
// C_AND/D//AND/D      x53y64     80'h00_FE00_80_0000_0C88_4F88
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a295_1 ( .OUT(na295_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1149_2), .IN8(na1718_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a295_2 ( .OUT(na295_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na295_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a295_4 ( .OUT(na295_2_i), .IN1(na221_1), .IN2(na295_1), .IN3(na297_2), .IN4(na4162_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a295_5 ( .OUT(na295_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na295_2_i) );
// C_AND/D//AND/D      x58y63     80'h00_FE00_80_0000_0C88_2F4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a297_1 ( .OUT(na297_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1720_1), .IN8(~na4366_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a297_2 ( .OUT(na297_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na297_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a297_4 ( .OUT(na297_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1149_2), .IN4(na1718_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a297_5 ( .OUT(na297_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na297_2_i) );
// C_MX4b/D///      x17y60     80'h00_FE00_00_0040_0A31_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a299_1 ( .OUT(na299_1_i), .IN1(~na310_2), .IN2(1'b1), .IN3(1'b1), .IN4(na214_2), .IN5(~na310_1), .IN6(na299_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a299_2 ( .OUT(na299_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na299_1_i) );
// C_ORAND////      x47y47     80'h00_0018_00_0000_0C88_3DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a301_1 ( .OUT(na301_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na266_1), .IN6(na4069_2), .IN7(1'b0), .IN8(~na302_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x44y48     80'h00_0018_00_0000_0C88_41FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a302_1 ( .OUT(na302_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na886_1), .IN6(~na122_1), .IN7(~na2529_2),
                     .IN8(na1495_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x18y54     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a303_4 ( .OUT(na303_2), .IN1(1'b1), .IN2(1'b1), .IN3(na952_2), .IN4(na4166_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x20y57     80'h00_0078_00_0000_0C88_548C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a304_1 ( .OUT(na304_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4528_2), .IN6(na2478_1), .IN7(~na2481_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a304_4 ( .OUT(na304_2), .IN1(1'b1), .IN2(na2478_2), .IN3(na2481_2), .IN4(na187_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x17y53     80'h00_0018_00_0040_0A17_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a307_1 ( .OUT(na307_1), .IN1(1'b1), .IN2(na4535_2), .IN3(~na4526_2), .IN4(1'b1), .IN5(~na3287_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x17y59     80'h00_0078_00_0000_0C88_322F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a310_1 ( .OUT(na310_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na307_1), .IN6(~na957_2), .IN7(1'b1), .IN8(~na303_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a310_4 ( .OUT(na310_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1567_1), .IN4(~na124_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x28y77     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a311_1 ( .OUT(na311_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na312_1), .IN6(na4167_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a311_2 ( .OUT(na311_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na311_1_i) );
// C_MX4b/D///      x27y77     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a312_1 ( .OUT(na312_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na312_1), .IN6(na313_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a312_2 ( .OUT(na312_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na312_1_i) );
// C_MX4b/D///      x29y78     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a313_1 ( .OUT(na313_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na314_1), .IN6(na313_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a313_2 ( .OUT(na313_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na313_1_i) );
// C_MX4b/D///      x29y77     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a314_1 ( .OUT(na314_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na314_1), .IN6(na1396_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a314_2 ( .OUT(na314_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na314_1_i) );
// C_MX4b/D///      x35y68     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a315_1 ( .OUT(na315_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na36_1), .IN6(na315_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a315_2 ( .OUT(na315_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na315_1_i) );
// C_MX4b/D///      x23y77     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a316_1 ( .OUT(na316_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na316_1), .IN6(na35_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a316_2 ( .OUT(na316_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na316_1_i) );
// C_///OR/      x22y67     80'h00_0060_00_0000_0C0E_FFCC
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a317_4 ( .OUT(na317_2), .IN1(1'b0), .IN2(na138_1), .IN3(1'b0), .IN4(na688_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x18y71     80'h00_0018_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a318_1 ( .OUT(na318_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na319_2), .IN8(~na4142_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y71     80'h00_0060_00_0000_0C08_FF51
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a319_4 ( .OUT(na319_2), .IN1(~na7_2), .IN2(~na2_1), .IN3(~na11_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x25y68     80'h00_0018_00_0000_0C88_ECFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a321_1 ( .OUT(na321_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na137_2), .IN7(na319_2), .IN8(na3292_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x36y72     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a322_1 ( .OUT(na322_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na323_1),
                     .IN8(na322_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a322_2 ( .OUT(na322_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na322_1_i) );
// C_MX4b/D///      x38y69     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a323_1 ( .OUT(na323_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na323_1), .IN8(na162_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a323_2 ( .OUT(na323_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na323_1_i) );
// C_MX4b/D///      x33y68     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a324_1 ( .OUT(na324_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na325_1), .IN6(na324_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a324_2 ( .OUT(na324_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na324_1_i) );
// C_MX4b/D///      x35y65     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a325_1 ( .OUT(na325_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na325_1), .IN6(na315_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a325_2 ( .OUT(na325_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na325_1_i) );
// C_ORAND*/D///      x50y63     80'h00_FE00_00_0000_0788_5FD3
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a326_1 ( .OUT(na326_1_i), .IN1(1'b0), .IN2(~na33_1), .IN3(~na326_1), .IN4(na4437_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na1149_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a326_2 ( .OUT(na326_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na326_1_i) );
// C_MX4b/D///      x52y78     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a327_1 ( .OUT(na327_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4169_2),
                     .IN8(na327_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a327_2 ( .OUT(na327_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na327_1_i) );
// C_MX4b/D///      x20y75     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a328_1 ( .OUT(na328_1_i), .IN1(1'b1), .IN2(na137_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na328_1),
                     .IN8(na3150_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a328_2 ( .OUT(na328_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na328_1_i) );
// C_MX4b/D///      x51y65     80'h00_FE00_00_0040_0A3C_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a329_1 ( .OUT(na329_1_i), .IN1(na1465_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na329_1), .IN6(na331_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a329_2 ( .OUT(na329_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na329_1_i) );
// C_MX4b/D///      x51y66     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a330_1 ( .OUT(na330_1_i), .IN1(~na1465_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na329_1), .IN6(na330_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a330_2 ( .OUT(na330_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na330_1_i) );
// C_MX4b/D///      x57y68     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a331_1 ( .OUT(na331_1_i), .IN1(~na1465_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na221_1), .IN6(na331_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a331_2 ( .OUT(na331_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na331_1_i) );
// C_MX4b/D///      x50y61     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a332_1 ( .OUT(na332_1_i), .IN1(~na1465_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na333_1), .IN6(na4172_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a332_2 ( .OUT(na332_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na332_1_i) );
// C_MX4b/D///      x45y59     80'h00_FE00_00_0040_0A32_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a333_1 ( .OUT(na333_1_i), .IN1(1'b1), .IN2(na346_2), .IN3(1'b1), .IN4(na4160_2), .IN5(na333_1), .IN6(~na346_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a333_2 ( .OUT(na333_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na333_1_i) );
// C_ORAND*////D      x51y61     80'h00_FE18_00_0000_0788_ADD3
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a335_1 ( .OUT(na335_1), .IN1(1'b0), .IN2(~na281_1), .IN3(~na790_2), .IN4(na336_2), .IN5(~na358_2), .IN6(na343_1), .IN7(na1570_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a335_5 ( .OUT(na335_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na335_1) );
// C_///ORAND/      x66y42     80'h00_0060_00_0000_0C08_FFD5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a336_4 ( .OUT(na336_2), .IN1(~na337_2), .IN2(1'b0), .IN3(~na80_1), .IN4(na338_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y39     80'h00_0060_00_0000_0C08_FF4A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a337_4 ( .OUT(na337_2), .IN1(na1473_2), .IN2(1'b1), .IN3(~na276_1), .IN4(na338_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y56     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a338_4 ( .OUT(na338_2), .IN1(~na709_1), .IN2(1'b1), .IN3(~na2278_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x52y64     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a340_4 ( .OUT(na340_2), .IN1(na785_2), .IN2(na341_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x59y60     80'h00_0078_00_0000_0C88_348A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a341_1 ( .OUT(na341_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2229_1), .IN6(na2228_2), .IN7(1'b1), .IN8(~na4511_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a341_4 ( .OUT(na341_2), .IN1(na2229_1), .IN2(1'b1), .IN3(na260_2), .IN4(na4511_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y62     80'h00_0018_00_0040_0A17_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a343_1 ( .OUT(na343_1), .IN1(1'b1), .IN2(~na2228_2), .IN3(1'b1), .IN4(na4510_2), .IN5(~na3298_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x51y64     80'h00_0078_00_0000_0C88_1C5A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a346_1 ( .OUT(na346_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na343_1), .IN7(~na790_2), .IN8(~na340_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a346_4 ( .OUT(na346_2), .IN1(na335_1), .IN2(1'b1), .IN3(~na332_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/D      x59y71     80'h00_FE00_80_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a349_4 ( .OUT(na349_2_i), .IN1(na350_1), .IN2(na3301_1), .IN3(~na1149_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a349_5 ( .OUT(na349_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na349_2_i) );
// C_MX4a////      x59y63     80'h00_0018_00_0040_0C14_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a350_1 ( .OUT(na350_1), .IN1(1'b1), .IN2(1'b0), .IN3(na3302_2), .IN4(1'b0), .IN5(1'b1), .IN6(~na357_1), .IN7(1'b1), .IN8(~na4511_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x71y55     80'h00_0018_00_0040_0CAA_1F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a351_1 ( .OUT(na351_1), .IN1(1'b0), .IN2(~na352_1), .IN3(1'b0), .IN4(~na4178_2), .IN5(1'b1), .IN6(1'b1), .IN7(~na2223_1),
                     .IN8(~na4504_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////D      x67y54     80'h00_FA18_00_0040_0AF1_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a352_1 ( .OUT(na352_1), .IN1(1'b1), .IN2(na4175_2), .IN3(1'b1), .IN4(na720_1), .IN5(~na355_1), .IN6(na1466_1), .IN7(na4433_2),
                     .IN8(na4177_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a352_5 ( .OUT(na352_2), .CLK(na1739_1), .EN(na1465_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na352_1) );
// C_MX2b////      x64y53     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a353_1 ( .OUT(na353_1), .IN1(1'b1), .IN2(~na2228_1), .IN3(1'b0), .IN4(1'b0), .IN5(na4176_2), .IN6(na3276_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x54y35     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a354_1 ( .OUT(na354_1), .IN1(1'b1), .IN2(~na273_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3726_1), .IN8(~na714_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x63y57     80'h00_0018_00_0000_0C88_DCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a355_1 ( .OUT(na355_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na295_2), .IN7(~na2223_1), .IN8(na3305_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x62y53     80'h00_0018_00_0000_0C88_6AFF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a356_1 ( .OUT(na356_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1465_1), .IN6(1'b0), .IN7(~na353_1), .IN8(na720_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x59y64     80'h00_0018_00_0000_0C88_48FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a357_1 ( .OUT(na357_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na333_1), .IN6(na295_2), .IN7(~na4507_2), .IN8(na4510_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x51y53     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a358_4 ( .OUT(na358_2_i), .IN1(na333_1), .IN2(na295_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a358_5 ( .OUT(na358_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na358_2_i) );
// C_AND/D//AND/D      x65y79     80'h00_FE00_80_0000_0C88_2F2F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a360_1 ( .OUT(na360_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1643_2), .IN8(~na4366_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a360_2 ( .OUT(na360_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na360_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a360_4 ( .OUT(na360_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1643_1), .IN4(~na4366_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a360_5 ( .OUT(na360_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na360_2_i) );
// C_MX4b/D///      x23y88     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a361_1 ( .OUT(na361_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na370_1), .IN6(na361_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a361_2 ( .OUT(na361_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na361_1_i) );
// C_MX2b////D      x58y67     80'h00_FA18_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a362_1 ( .OUT(na362_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4153_2), .IN5(na543_1), .IN6(1'b0), .IN7(na3151_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a362_5 ( .OUT(na362_2), .CLK(na1739_1), .EN(na372_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na362_1) );
// C_MX2b////D      x54y65     80'h00_FA18_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a363_1 ( .OUT(na363_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4153_2), .IN5(na543_2), .IN6(1'b0), .IN7(na3152_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a363_5 ( .OUT(na363_2), .CLK(na1739_1), .EN(na372_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na363_1) );
// C_MX2b////D      x50y68     80'h00_FA18_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a364_1 ( .OUT(na364_1), .IN1(1'b1), .IN2(~na285_1), .IN3(1'b0), .IN4(1'b0), .IN5(na545_1), .IN6(na3153_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a364_5 ( .OUT(na364_2), .CLK(na1739_1), .EN(na372_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na364_1) );
// C_MX2b////D      x54y69     80'h00_FA18_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a365_1 ( .OUT(na365_1), .IN1(1'b1), .IN2(~na285_1), .IN3(1'b0), .IN4(1'b0), .IN5(na545_2), .IN6(na3154_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a365_5 ( .OUT(na365_2), .CLK(na1739_1), .EN(na372_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na365_1) );
// C_MX2b////D      x56y68     80'h00_FA18_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a366_1 ( .OUT(na366_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4153_2), .IN5(na3155_1), .IN6(1'b0), .IN7(na547_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a366_5 ( .OUT(na366_2), .CLK(na1739_1), .EN(na372_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na366_1) );
// C_MX2b////D      x52y63     80'h00_FA18_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a367_1 ( .OUT(na367_1), .IN1(1'b1), .IN2(~na285_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na547_2), .IN8(na3156_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a367_5 ( .OUT(na367_2), .CLK(na1739_1), .EN(na372_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na367_1) );
// C_MX2b////D      x54y67     80'h00_FA18_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a368_1 ( .OUT(na368_1), .IN1(1'b1), .IN2(~na285_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na549_1), .IN8(na3157_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a368_5 ( .OUT(na368_2), .CLK(na1739_1), .EN(na372_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na368_1) );
// C_MX2b////D      x56y70     80'h00_FA18_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a369_1 ( .OUT(na369_1), .IN1(1'b1), .IN2(~na285_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na549_2), .IN8(na3158_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a369_5 ( .OUT(na369_2), .CLK(na1739_1), .EN(na372_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na369_1) );
// C_MX4b/D///      x23y89     80'h00_FE00_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a370_1 ( .OUT(na370_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4189_2),
                     .IN8(na371_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a370_2 ( .OUT(na370_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na370_1_i) );
// C_MX4b/D///      x26y88     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a371_1 ( .OUT(na371_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na4190_2), .IN6(na373_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a371_2 ( .OUT(na371_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na371_1_i) );
// C_AND////      x49y75     80'h00_0018_00_0000_0C88_4AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a372_1 ( .OUT(na372_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4400_2), .IN6(1'b1), .IN7(~na287_2), .IN8(na1296_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x23y90     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a373_1 ( .OUT(na373_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na374_1), .IN6(na373_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a373_2 ( .OUT(na373_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na373_1_i) );
// C_MX4b/D///      x21y89     80'h00_FE00_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a374_1 ( .OUT(na374_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na384_1),
                     .IN8(na4191_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a374_2 ( .OUT(na374_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na374_1_i) );
// C_MX2b/D///      x43y77     80'h00_F600_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a375_1 ( .OUT(na375_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na376_1), .IN5(na4181_2), .IN6(1'b0), .IN7(na362_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a375_2 ( .OUT(na375_1), .CLK(na1739_1), .EN(~na1398_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na375_1_i) );
// C_ORAND////      x38y76     80'h00_0018_00_0000_0C88_BAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a376_1 ( .OUT(na376_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4400_2), .IN6(1'b0), .IN7(na287_2), .IN8(~na1296_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x42y75     80'h00_F600_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a377_1 ( .OUT(na377_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na376_1), .IN5(na4182_2), .IN6(1'b0), .IN7(na363_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a377_2 ( .OUT(na377_1), .CLK(na1739_1), .EN(~na1398_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na377_1_i) );
// C_MX2b/D///      x37y72     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a378_1 ( .OUT(na378_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na376_1), .IN5(1'b0), .IN6(na4183_2), .IN7(1'b0), .IN8(na364_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a378_2 ( .OUT(na378_1), .CLK(na1739_1), .EN(~na1398_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na378_1_i) );
// C_MX2b/D///      x41y73     80'h00_F600_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a379_1 ( .OUT(na379_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na376_1), .IN5(na4184_2), .IN6(1'b0), .IN7(na365_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a379_2 ( .OUT(na379_1), .CLK(na1739_1), .EN(~na1398_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na379_1_i) );
// C_MX2b/D///      x44y74     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a380_1 ( .OUT(na380_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na376_1), .IN5(1'b0), .IN6(na4185_2), .IN7(1'b0), .IN8(na366_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a380_2 ( .OUT(na380_1), .CLK(na1739_1), .EN(~na1398_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na380_1_i) );
// C_MX2b/D///      x42y73     80'h00_F600_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a381_1 ( .OUT(na381_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na376_1), .IN5(na4186_2), .IN6(1'b0), .IN7(na367_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a381_2 ( .OUT(na381_1), .CLK(na1739_1), .EN(~na1398_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na381_1_i) );
// C_MX2b/D///      x43y76     80'h00_F600_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a382_1 ( .OUT(na382_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na376_1), .IN5(na4187_2), .IN6(1'b0), .IN7(na368_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a382_2 ( .OUT(na382_1), .CLK(na1739_1), .EN(~na1398_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na382_1_i) );
// C_MX2b/D///      x42y78     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a383_1 ( .OUT(na383_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na376_1), .IN5(1'b0), .IN6(na4188_2), .IN7(1'b0), .IN8(na369_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a383_2 ( .OUT(na383_1), .CLK(na1739_1), .EN(~na1398_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na383_1_i) );
// C_MX4b/D///      x24y91     80'h00_FE00_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a384_1 ( .OUT(na384_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na384_1),
                     .IN8(na1332_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a384_2 ( .OUT(na384_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na384_1_i) );
// C_///AND/D      x13y84     80'h00_FE00_80_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a387_4 ( .OUT(na387_2_i), .IN1(na1666_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1347_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a387_5 ( .OUT(na387_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na387_2_i) );
// C_AND/D//AND/D      x18y89     80'h00_FE00_80_0000_0C88_3A1F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a388_1 ( .OUT(na388_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1666_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1347_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a388_2 ( .OUT(na388_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na388_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a388_4 ( .OUT(na388_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na388_2), .IN4(~na1347_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a388_5 ( .OUT(na388_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na388_2_i) );
// C_AND/D//AND/D      x19y89     80'h00_FE00_80_0000_0C88_3C3C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a390_1 ( .OUT(na390_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1668_2), .IN7(1'b1), .IN8(~na1347_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a390_2 ( .OUT(na390_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na390_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a390_4 ( .OUT(na390_2_i), .IN1(1'b1), .IN2(na1668_1), .IN3(1'b1), .IN4(~na1347_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a390_5 ( .OUT(na390_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na390_2_i) );
// C_AND/D//ORAND*/D      x25y92     80'h00_FE00_80_0000_0C87_3AD3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a391_1 ( .OUT(na391_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1670_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1347_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a391_2 ( .OUT(na391_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na391_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a391_4 ( .OUT(na391_2_i), .IN1(1'b0), .IN2(~na391_1), .IN3(~na1511_2), .IN4(na2707_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a391_5 ( .OUT(na391_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na391_2_i) );
// C_AND/D///      x50y78     80'h00_FE00_00_0000_0888_1221
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a392_1 ( .OUT(na392_1_i), .IN1(~na456_1), .IN2(~na4367_2), .IN3(na9_1), .IN4(~na392_1), .IN5(na145_1), .IN6(~na285_1), .IN7(~na9_2),
                     .IN8(~na4154_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a392_2 ( .OUT(na392_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na392_1_i) );
// C_ORAND////      x15y65     80'h00_0018_00_0000_0C88_AEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a394_1 ( .OUT(na394_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1614_1), .IN6(na405_2), .IN7(na4474_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x14y65     80'h00_0060_00_0000_0C08_FFCE
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a395_4 ( .OUT(na395_2), .IN1(na4470_2), .IN2(na2_2), .IN3(1'b0), .IN4(na1610_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x22y72     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a396_1 ( .OUT(na396_1_i), .IN1(1'b1), .IN2(~na137_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3160_1),
                     .IN8(na396_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a396_2 ( .OUT(na396_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na396_1_i) );
// C_AND/D///      x40y55     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a397_1 ( .OUT(na397_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na399_2), .IN6(1'b1), .IN7(1'b1), .IN8(na3413_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a397_2 ( .OUT(na397_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na397_1_i) );
// C_AND/D///      x42y55     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a398_1 ( .OUT(na398_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na399_1), .IN6(1'b1), .IN7(1'b1), .IN8(na3413_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a398_2 ( .OUT(na398_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na398_1_i) );
// C_AND////D      x41y61     80'h00_FE18_00_0000_0888_F35C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a399_1 ( .OUT(na399_1), .IN1(1'b1), .IN2(na403_2), .IN3(~na402_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na403_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a399_5 ( .OUT(na399_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na399_1) );
// C_///AND/D      x52y83     80'h00_FE00_80_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a402_4 ( .OUT(na402_2_i), .IN1(~na218_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1678_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a402_5 ( .OUT(na402_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na402_2_i) );
// C_AND/D//AND/D      x45y82     80'h00_FE00_80_0000_0C88_C5F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a403_1 ( .OUT(na403_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na218_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1678_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a403_2 ( .OUT(na403_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na403_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a403_4 ( .OUT(na403_2_i), .IN1(~na218_1), .IN2(~na403_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a403_5 ( .OUT(na403_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na403_2_i) );
// C_///ORAND/      x25y68     80'h00_0060_00_0000_0C08_FFE3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a405_4 ( .OUT(na405_2), .IN1(1'b0), .IN2(~na138_1), .IN3(na407_2), .IN4(na3310_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x34y63     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a407_4 ( .OUT(na407_2), .IN1(~na1290_1), .IN2(1'b1), .IN3(na8_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y71     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a408_1 ( .OUT(na408_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na984_1), .IN6(na12_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x50y90     80'h00_FE00_00_0040_0AC8_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a409_1 ( .OUT(na409_1_i), .IN1(na430_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4192_2),
                     .IN8(~na409_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a409_2 ( .OUT(na409_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na409_1_i) );
// C_MX4b/D///      x41y87     80'h00_FE00_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a410_1 ( .OUT(na410_1_i), .IN1(~na430_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1685_1),
                     .IN8(na4193_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a410_2 ( .OUT(na410_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na410_1_i) );
// C_MX2b/D///      x17y85     80'h00_F600_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a411_1 ( .OUT(na411_1_i), .IN1(1'b1), .IN2(na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na375_1), .IN6(na412_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a411_2 ( .OUT(na411_1), .CLK(na1739_1), .EN(~na1418_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na411_1_i) );
// C_MX2b/D///      x21y82     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a412_1 ( .OUT(na412_1_i), .IN1(1'b1), .IN2(na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na377_1), .IN8(na413_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a412_2 ( .OUT(na412_1), .CLK(na1739_1), .EN(~na1418_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na412_1_i) );
// C_MX2b/D///      x22y80     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a413_1 ( .OUT(na413_1_i), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na414_1), .IN6(na378_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a413_2 ( .OUT(na413_1), .CLK(na1739_1), .EN(~na1418_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na413_1_i) );
// C_MX2b/D///      x25y79     80'h00_F600_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a414_1 ( .OUT(na414_1_i), .IN1(1'b1), .IN2(na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na379_1), .IN6(na415_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a414_2 ( .OUT(na414_1), .CLK(na1739_1), .EN(~na1418_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na414_1_i) );
// C_MX2b/D///      x25y78     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a415_1 ( .OUT(na415_1_i), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na416_1), .IN8(na380_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a415_2 ( .OUT(na415_1), .CLK(na1739_1), .EN(~na1418_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na415_1_i) );
// C_MX2b/D///      x26y79     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a416_1 ( .OUT(na416_1_i), .IN1(1'b1), .IN2(na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na381_1), .IN8(na417_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a416_2 ( .OUT(na416_1), .CLK(na1739_1), .EN(~na1418_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na416_1_i) );
// C_MX2b/D///      x26y82     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a417_1 ( .OUT(na417_1_i), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(na418_1), .IN6(na382_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a417_2 ( .OUT(na417_1), .CLK(na1739_1), .EN(~na1418_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na417_1_i) );
// C_MX2b/D///      x21y83     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a418_1 ( .OUT(na418_1_i), .IN1(1'b1), .IN2(~na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1351_2), .IN8(na383_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a418_2 ( .OUT(na418_1), .CLK(na1739_1), .EN(~na1418_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na418_1_i) );
// C_///AND/      x28y70     80'h00_0060_00_0000_0C08_FF51
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a420_4 ( .OUT(na420_2), .IN1(~na7_2), .IN2(~na2_1), .IN3(~na3312_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x23y64     80'h00_0018_00_0000_0888_FE3C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a421_1 ( .OUT(na421_1), .IN1(1'b0), .IN2(na3313_1), .IN3(1'b0), .IN4(~na1539_1), .IN5(na425_2), .IN6(na423_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x25y66     80'h00_0078_00_0000_0C88_A3F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a423_1 ( .OUT(na423_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na424_2), .IN7(na531_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a423_4 ( .OUT(na423_2), .IN1(~na425_2), .IN2(~na423_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x33y82     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a424_4 ( .OUT(na424_2), .IN1(na456_1), .IN2(1'b1), .IN3(~na443_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x51y81     80'h00_0060_00_0000_0C08_FF21
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a425_4 ( .OUT(na425_2), .IN1(~na456_1), .IN2(~na4372_2), .IN3(na9_1), .IN4(~na3014_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x32y67     80'h00_FE00_00_0000_0C88_2CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a426_1 ( .OUT(na426_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na929_1), .IN7(na928_1), .IN8(~na926_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a426_2 ( .OUT(na426_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na426_1_i) );
// C_OR////D      x25y56     80'h00_FE18_00_0000_0EEE_03C0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a427_1 ( .OUT(na427_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3316_1), .IN5(1'b0), .IN6(~na421_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a427_5 ( .OUT(na427_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na427_1) );
// C_MX4b/D///      x57y74     80'h00_FE00_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a428_1 ( .OUT(na428_1_i), .IN1(~na105_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1630_1),
                     .IN8(na4196_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a428_2 ( .OUT(na428_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na428_1_i) );
// C_MX4b/D///      x44y88     80'h00_FE00_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a429_1 ( .OUT(na429_1_i), .IN1(~na430_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1685_2),
                     .IN8(na429_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a429_2 ( .OUT(na429_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na429_1_i) );
// C_///ORAND/D      x47y89     80'h00_FE00_80_0000_0C08_FFAE
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a430_4 ( .OUT(na430_2_i), .IN1(na430_2), .IN2(na4138_2), .IN3(na3317_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a430_5 ( .OUT(na430_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na430_2_i) );
// C_///AND/D      x36y87     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a432_4 ( .OUT(na432_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1149_2), .IN4(na1674_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a432_5 ( .OUT(na432_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na432_2_i) );
// C_AND/D//AND/D      x35y91     80'h00_FE00_80_0000_0C88_2F4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a434_1 ( .OUT(na434_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1676_1), .IN8(~na4366_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a434_2 ( .OUT(na434_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na434_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a434_4 ( .OUT(na434_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1149_2), .IN4(na1674_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a434_5 ( .OUT(na434_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na434_2_i) );
// C_AND/D//AND/D      x35y73     80'h00_FE00_80_0000_0C88_5A5A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a435_1 ( .OUT(na435_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na436_1), .IN6(1'b1), .IN7(~na1149_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a435_2 ( .OUT(na435_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na435_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a435_4 ( .OUT(na435_2_i), .IN1(na435_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a435_5 ( .OUT(na435_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na435_2_i) );
// C_AND////      x33y65     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a436_1 ( .OUT(na436_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na423_1), .IN7(1'b1), .IN8(na1539_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x48y42     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a437_1 ( .OUT(na437_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4228_2), .IN5(na438_1), .IN6(1'b0), .IN7(na3717_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a437_2 ( .OUT(na437_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na437_1_i) );
// C_MX2b/D///      x49y39     80'h00_FE00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a438_1 ( .OUT(na438_1_i), .IN1(1'b1), .IN2(na536_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na439_1), .IN8(na3716_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a438_2 ( .OUT(na438_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na438_1_i) );
// C_MX2b/D///      x50y39     80'h00_FE00_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a439_1 ( .OUT(na439_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4228_2), .IN5(1'b0), .IN6(na440_1), .IN7(1'b0), .IN8(na3715_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a439_2 ( .OUT(na439_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na439_1_i) );
// C_MX2b/D///      x47y40     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a440_1 ( .OUT(na440_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4228_2), .IN5(na441_1), .IN6(1'b0), .IN7(na3714_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a440_2 ( .OUT(na440_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na440_1_i) );
// C_MX2b/D///      x47y37     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a441_1 ( .OUT(na441_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4228_2), .IN5(na442_1), .IN6(1'b0), .IN7(na3713_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a441_2 ( .OUT(na441_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na441_1_i) );
// C_MX2b/D///      x45y39     80'h00_FE00_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a442_1 ( .OUT(na442_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4228_2), .IN5(1'b0), .IN6(na84_2), .IN7(1'b0), .IN8(na3712_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a442_2 ( .OUT(na442_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na442_1_i) );
// C_MX4b/D///      x62y89     80'h00_FE00_00_0040_0A51_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a443_1 ( .OUT(na443_1_i), .IN1(na456_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4204_2), .IN5(~na455_1), .IN6(1'b0), .IN7(na443_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a443_2 ( .OUT(na443_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na443_1_i) );
// C_ORAND*////D      x51y83     80'h00_FE18_00_0000_0788_ABB5
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a445_1 ( .OUT(na445_1), .IN1(~na435_2), .IN2(1'b0), .IN3(na446_2), .IN4(~na4398_2), .IN5(na452_1), .IN6(~na469_2), .IN7(na1574_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a445_5 ( .OUT(na445_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na445_1) );
// C_///ORAND/      x40y63     80'h00_0060_00_0000_0C08_FFB5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a446_4 ( .OUT(na446_2), .IN1(~na447_2), .IN2(1'b0), .IN3(na9_2), .IN4(~na392_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y61     80'h00_0060_00_0000_0C08_FF12
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a447_4 ( .OUT(na447_2), .IN1(na4460_2), .IN2(~na423_1), .IN3(~na1198_1), .IN4(~na3014_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y83     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a449_4 ( .OUT(na449_2), .IN1(na1255_2), .IN2(1'b1), .IN3(1'b1), .IN4(na450_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x56y88     80'h00_0078_00_0000_0C88_32A8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a450_1 ( .OUT(na450_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2962_1), .IN6(~na2965_2), .IN7(1'b1), .IN8(~na4571_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a450_4 ( .OUT(na450_2), .IN1(na2962_2), .IN2(na2965_2), .IN3(na1269_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y87     80'h00_0018_00_0040_0A4D_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a452_1 ( .OUT(na452_1), .IN1(1'b1), .IN2(na2965_2), .IN3(1'b1), .IN4(na4568_2), .IN5(1'b1), .IN6(1'b0), .IN7(~na3324_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x57y89     80'h00_0078_00_0000_0C88_523C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a455_1 ( .OUT(na455_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na452_1), .IN6(~na1260_2), .IN7(~na449_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a455_4 ( .OUT(na455_2), .IN1(1'b1), .IN2(na4203_2), .IN3(1'b1), .IN4(~na518_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D//AND/D      x53y77     80'h00_FE00_80_0000_0C88_5E88
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a456_1 ( .OUT(na456_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na456_1), .IN6(na4202_2), .IN7(~na4206_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a456_2 ( .OUT(na456_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na456_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a456_4 ( .OUT(na456_2_i), .IN1(na507_1), .IN2(na4333_2), .IN3(na980_2), .IN4(na986_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a456_5 ( .OUT(na456_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na456_2_i) );
// C_ORAND/D///      x49y87     80'h00_FE00_00_0000_0C88_5EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a457_1 ( .OUT(na457_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na458_1), .IN6(na3327_1), .IN7(~na1149_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a457_2 ( .OUT(na457_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na457_1_i) );
// C_MX4a////      x59y89     80'h00_0018_00_0040_0C28_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a458_1 ( .OUT(na458_1), .IN1(1'b0), .IN2(1'b1), .IN3(1'b0), .IN4(na3328_2), .IN5(1'b1), .IN6(na468_2), .IN7(1'b1), .IN8(~na4571_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x66y85     80'h00_0018_00_0040_0C55_1000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a459_1 ( .OUT(na459_1), .IN1(~na460_1), .IN2(1'b0), .IN3(~na467_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na2958_2),
                     .IN8(~na4565_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////D      x65y85     80'h00_FA18_00_0040_0AF4_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a460_1 ( .OUT(na460_1), .IN1(1'b1), .IN2(na4209_2), .IN3(1'b1), .IN4(~na1388_1), .IN5(na1532_1), .IN6(na466_1), .IN7(~na4211_2),
                     .IN8(na4456_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a460_5 ( .OUT(na460_2), .CLK(na1739_1), .EN(na456_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na460_1) );
// C_MX2b////      x66y83     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a461_1 ( .OUT(na461_1), .IN1(~na2963_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na465_1), .IN8(na3329_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x56y83     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a462_1 ( .OUT(na462_1), .IN1(na463_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4207_2), .IN5(na1156_1), .IN6(na1151_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x59y85     80'h00_0018_00_0000_0C88_12FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a463_1 ( .OUT(na463_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2963_2), .IN6(~na4569_2), .IN7(~na2961_1),
                     .IN8(~na4568_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x38y55     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a465_1 ( .OUT(na465_1), .IN1(~na888_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3444_1), .IN8(~na1358_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x63y84     80'h00_0018_00_0000_0C88_DAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a466_1 ( .OUT(na466_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na456_2), .IN6(1'b0), .IN7(~na2958_1), .IN8(na3331_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x68y83     80'h00_0018_00_0000_0C88_6AFF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a467_1 ( .OUT(na467_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1531_2), .IN6(1'b0), .IN7(~na461_1), .IN8(na1388_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y84     80'h00_0060_00_0000_0C08_FF28
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a468_4 ( .OUT(na468_2), .IN1(na456_2), .IN2(na2965_2), .IN3(na443_1), .IN4(~na4568_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x51y86     80'h00_FE00_80_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a469_4 ( .OUT(na469_2_i), .IN1(na456_2), .IN2(1'b1), .IN3(na443_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a469_5 ( .OUT(na469_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na469_2_i) );
// C_MX2b/D///      x63y64     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a470_1 ( .OUT(na470_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2124_1), .IN8(na471_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a470_2 ( .OUT(na470_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na470_1_i) );
// C_MX2b/D///      x60y62     80'h00_F600_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a471_1 ( .OUT(na471_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1887_2), .IN6(na472_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a471_2 ( .OUT(na471_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na471_1_i) );
// C_MX2b/D///      x61y58     80'h00_F600_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a472_1 ( .OUT(na472_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1443_2), .IN5(na1887_1), .IN6(1'b0), .IN7(na473_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a472_2 ( .OUT(na472_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na472_1_i) );
// C_MX2b/D///      x60y57     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a473_1 ( .OUT(na473_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1443_2), .IN5(na474_1), .IN6(1'b0), .IN7(na1889_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a473_2 ( .OUT(na473_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na473_1_i) );
// C_MX2b/D///      x55y57     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a474_1 ( .OUT(na474_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1889_1), .IN8(na480_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a474_2 ( .OUT(na474_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na474_1_i) );
// C_MX2b/D///      x67y63     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a475_1 ( .OUT(na475_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1866_2), .IN8(na476_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a475_2 ( .OUT(na475_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na475_1_i) );
// C_MX2b/D///      x62y64     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a476_1 ( .OUT(na476_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1443_2), .IN5(na477_1), .IN6(1'b0), .IN7(na1866_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a476_2 ( .OUT(na476_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na476_1_i) );
// C_MX2b/D///      x59y57     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a477_1 ( .OUT(na477_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1868_2), .IN8(na478_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a477_2 ( .OUT(na477_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na477_1_i) );
// C_MX2b/D///      x56y58     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a478_1 ( .OUT(na478_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1868_1), .IN8(na479_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a478_2 ( .OUT(na478_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na478_1_i) );
// C_MX2b/D///      x48y50     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a479_1 ( .OUT(na479_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3718_1), .IN8(na480_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a479_2 ( .OUT(na479_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na479_1_i) );
// C_MX2b/D///      x50y50     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a480_1 ( .OUT(na480_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1443_2), .IN5(na481_1), .IN6(1'b0), .IN7(na3717_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a480_2 ( .OUT(na480_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na480_1_i) );
// C_MX2b/D///      x51y47     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a481_1 ( .OUT(na481_1_i), .IN1(1'b1), .IN2(~na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na482_1), .IN8(na3716_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a481_2 ( .OUT(na481_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na481_1_i) );
// C_MX2b/D///      x50y47     80'h00_F600_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a482_1 ( .OUT(na482_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1443_2), .IN5(1'b0), .IN6(na483_1), .IN7(1'b0), .IN8(na3715_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a482_2 ( .OUT(na482_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na482_1_i) );
// C_MX2b/D///      x49y48     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a483_1 ( .OUT(na483_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3714_1), .IN8(na484_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a483_2 ( .OUT(na483_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na483_1_i) );
// C_MX2b/D///      x50y48     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a484_1 ( .OUT(na484_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1443_2), .IN5(na1579_1), .IN6(1'b0), .IN7(na3713_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a484_2 ( .OUT(na484_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na484_1_i) );
// C_MX2b/D///      x64y64     80'h00_F600_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a485_1 ( .OUT(na485_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b0), .IN4(1'b0), .IN5(na4502_2), .IN6(na1993_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a485_2 ( .OUT(na485_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na485_1_i) );
// C_MX2b/D///      x69y63     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a486_1 ( .OUT(na486_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1866_2), .IN8(na487_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a486_2 ( .OUT(na486_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na486_1_i) );
// C_MX2b/D///      x68y62     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a487_1 ( .OUT(na487_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1891_2), .IN8(na488_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a487_2 ( .OUT(na487_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na487_1_i) );
// C_MX2b/D///      x66y62     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a488_1 ( .OUT(na488_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1443_2), .IN5(na489_1), .IN6(1'b0), .IN7(na1891_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a488_2 ( .OUT(na488_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na488_1_i) );
// C_MX2b/D///      x65y61     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a489_1 ( .OUT(na489_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1443_2), .IN5(na490_1), .IN6(1'b0), .IN7(na1893_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a489_2 ( .OUT(na489_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na489_1_i) );
// C_MX2b/D///      x65y59     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a490_1 ( .OUT(na490_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1443_2), .IN5(na491_1), .IN6(1'b0), .IN7(na1893_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a490_2 ( .OUT(na490_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na490_1_i) );
// C_MX2b/D///      x67y59     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a491_1 ( .OUT(na491_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1443_2), .IN5(na492_1), .IN6(1'b0), .IN7(na1862_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a491_2 ( .OUT(na491_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na491_1_i) );
// C_MX2b/D///      x63y59     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a492_1 ( .OUT(na492_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1443_2), .IN5(na493_1), .IN6(1'b0), .IN7(na1862_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a492_2 ( .OUT(na492_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na492_1_i) );
// C_MX2b/D///      x61y61     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a493_1 ( .OUT(na493_1_i), .IN1(1'b1), .IN2(na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1864_2), .IN8(na494_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a493_2 ( .OUT(na493_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na493_1_i) );
// C_MX2b/D///      x66y60     80'h00_F600_00_0040_0A51_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a494_1 ( .OUT(na494_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1443_2), .IN5(~na495_1), .IN6(1'b0), .IN7(na1864_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a494_2 ( .OUT(na494_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na494_1_i) );
// C_MX2b////      x63y67     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a495_1 ( .OUT(na495_1), .IN1(1'b1), .IN2(na1993_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na475_1), .IN6(~na1993_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x67y61     80'h00_FE00_00_0040_0A54_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a496_1 ( .OUT(na496_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na498_1), .IN5(na499_1), .IN6(1'b0), .IN7(~na497_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a496_2 ( .OUT(na496_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na496_1_i) );
// C_MX2b////      x70y57     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a497_1 ( .OUT(na497_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na54_2), .IN5(~na496_1), .IN6(1'b0), .IN7(~na1893_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x68y64     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a498_1 ( .OUT(na498_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4423_2), .IN6(na1986_2), .IN7(na4493_2), .IN8(na1990_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x69y57     80'h00_FE00_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a499_1 ( .OUT(na499_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na498_1), .IN5(na501_1), .IN6(1'b0), .IN7(na500_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a499_2 ( .OUT(na499_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na499_1_i) );
// C_MX2b////      x66y55     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a500_1 ( .OUT(na500_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na54_2), .IN5(na499_1), .IN6(1'b0), .IN7(na1862_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x69y59     80'h00_FE00_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a501_1 ( .OUT(na501_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na498_1), .IN5(na503_1), .IN6(1'b0), .IN7(na502_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a501_2 ( .OUT(na501_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na501_1_i) );
// C_MX2b////      x64y55     80'h00_0018_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a502_1 ( .OUT(na502_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na54_2), .IN5(na501_1), .IN6(1'b0), .IN7(na1862_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x63y61     80'h00_FE00_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a503_1 ( .OUT(na503_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na498_1), .IN5(na505_1), .IN6(1'b0), .IN7(na504_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a503_2 ( .OUT(na503_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na503_1_i) );
// C_MX2a////      x64y57     80'h00_0018_00_0040_0C05_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a504_1 ( .OUT(na504_1), .IN1(na503_1), .IN2(1'b0), .IN3(na1864_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na54_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x65y57     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a505_1 ( .OUT(na505_1_i), .IN1(na4084_2), .IN2(1'b1), .IN3(1'b1), .IN4(na498_1), .IN5(na505_1), .IN6(na4480_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a505_2 ( .OUT(na505_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na505_1_i) );
// C_///ORAND/D      x46y79     80'h00_FE00_80_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a506_4 ( .OUT(na506_2_i), .IN1(na4110_2), .IN2(~na138_1), .IN3(~na1149_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a506_5 ( .OUT(na506_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na506_2_i) );
// C_MX4b/D///      x53y85     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a507_1 ( .OUT(na507_1_i), .IN1(na456_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na507_1), .IN6(na1321_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a507_2 ( .OUT(na507_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na507_1_i) );
// C_///ORAND/D      x37y70     80'h00_FE00_80_0000_0C08_FF5D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a508_4 ( .OUT(na508_2_i), .IN1(~na3334_1), .IN2(na3335_1), .IN3(~na1149_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a508_5 ( .OUT(na508_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na508_2_i) );
// C_MX4b/D///      x53y90     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a510_1 ( .OUT(na510_1_i), .IN1(~na456_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na507_1), .IN6(na510_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a510_2 ( .OUT(na510_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na510_1_i) );
// C_MX4b////D      x68y69     80'h00_FA18_00_0040_0AF1_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a511_1 ( .OUT(na511_1), .IN1(1'b1), .IN2(na512_1), .IN3(na4226_2), .IN4(1'b1), .IN5(~na4218_2), .IN6(na4425_2), .IN7(na1444_1),
                     .IN8(na517_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a511_5 ( .OUT(na511_2), .CLK(na1739_1), .EN(na1443_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na511_1) );
// C_MX2b////      x67y72     80'h00_0018_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a512_1 ( .OUT(na512_1), .IN1(1'b1), .IN2(1'b1), .IN3(na1991_1), .IN4(1'b1), .IN5(1'b0), .IN6(na3336_1), .IN7(1'b0), .IN8(na4217_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x61y69     80'h00_0018_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a513_1 ( .OUT(na513_1), .IN1(na514_2), .IN2(1'b1), .IN3(na38_2), .IN4(1'b1), .IN5(na475_1), .IN6(na470_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y69     80'h00_0060_00_0000_0C08_FF21
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a514_4 ( .OUT(na514_2), .IN1(~na4489_2), .IN2(~na1989_2), .IN3(na1991_1), .IN4(~na1990_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x53y45     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a516_1 ( .OUT(na516_1), .IN1(1'b1), .IN2(~na536_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3718_1), .IN8(~na437_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x68y78     80'h00_0060_00_0000_0C08_FFAB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a517_4 ( .OUT(na517_2), .IN1(na3338_2), .IN2(~na1986_1), .IN3(na38_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x58y88     80'h00_FE00_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a518_1 ( .OUT(na518_1_i), .IN1(~na456_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na443_1),
                     .IN8(na518_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a518_2 ( .OUT(na518_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na518_1_i) );
// C_ANDXOR////D      x70y68     80'h00_FA18_00_0000_0666_F35D
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a519_1 ( .OUT(na519_1), .IN1(na535_1), .IN2(~na3341_1), .IN3(na520_2), .IN4(1'b1), .IN5(1'b1), .IN6(na1438_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a519_5 ( .OUT(na519_2), .CLK(na1739_1), .EN(na1436_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na519_1) );
// C_///AND/      x70y75     80'h00_0060_00_0000_0C08_FF13
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a520_4 ( .OUT(na520_2), .IN1(1'b1), .IN2(~na3336_1), .IN3(~na521_1), .IN4(~na1990_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x70y73     80'h00_0018_00_0000_0888_9FAC
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a521_1 ( .OUT(na521_1), .IN1(1'b0), .IN2(~na1993_2), .IN3(~na4221_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na4487_2),
                     .IN8(na1990_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x71y77     80'h00_0060_00_0000_0C08_FFC4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a522_4 ( .OUT(na522_2), .IN1(~na360_2), .IN2(na103_1), .IN3(1'b1), .IN4(na4222_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x65y80     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a523_1 ( .OUT(na523_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na360_1), .IN6(1'b1), .IN7(~na38_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x65y69     80'h00_0018_00_0000_0C88_ABFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a524_1 ( .OUT(na524_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3342_2), .IN6(~na1993_2), .IN7(na4226_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x63y71     80'h00_F600_00_0040_0C0C_F200
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a525_1 ( .OUT(na525_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na4219_2), .IN4(na2011_1), .IN5(na95_1), .IN6(~na4102_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a525_2 ( .OUT(na525_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na525_1_i) );
// C_ORAND////      x54y54     80'h00_0018_00_0000_0888_EFA3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a526_1 ( .OUT(na526_1), .IN1(1'b0), .IN2(~na1451_1), .IN3(na3343_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na528_1), .IN8(na55_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y61     80'h00_0018_00_0000_0C88_2CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a528_1 ( .OUT(na528_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na22_1), .IN7(na93_1), .IN8(~na1443_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x68y57     80'h00_FE00_80_0000_0C08_FF2A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a529_4 ( .OUT(na529_2_i), .IN1(na109_1), .IN2(1'b1), .IN3(na107_1), .IN4(~na104_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a529_5 ( .OUT(na529_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na529_2_i) );
// C_OR////D      x46y43     80'h00_FE18_00_0000_0EEE_B000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a530_1 ( .OUT(na530_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3346_1), .IN8(~na526_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a530_5 ( .OUT(na530_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na530_1) );
// C_ORAND*/D///      x36y75     80'h00_FE00_00_0000_0788_5FD3
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a531_1 ( .OUT(na531_1_i), .IN1(1'b0), .IN2(~na424_2), .IN3(~na531_1), .IN4(na1539_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1149_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a531_2 ( .OUT(na531_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na531_1_i) );
// C_MX4b/D///      x40y88     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a532_1 ( .OUT(na532_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4225_2),
                     .IN8(na532_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a532_2 ( .OUT(na532_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na532_1_i) );
// C_MX4b/D///      x29y81     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a533_1 ( .OUT(na533_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na533_1), .IN6(na1320_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a533_2 ( .OUT(na533_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na533_1_i) );
// C_ANDXOR/D//AND/D      x69y79     80'h00_FA00_80_0000_0C68_CEFA
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a534_1 ( .OUT(na534_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na4590_2), .IN6(~na1986_2), .IN7(1'b1), .IN8(~na4216_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a534_2 ( .OUT(na534_1), .CLK(na1739_1), .EN(na1435_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na534_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a534_4 ( .OUT(na534_2_i), .IN1(na534_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a534_5 ( .OUT(na534_2), .CLK(na1739_1), .EN(na1435_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na534_2_i) );
// C_MX2b/D///      x65y63     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a535_1 ( .OUT(na535_1_i), .IN1(1'b1), .IN2(~na536_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3718_1), .IN8(na537_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a535_2 ( .OUT(na535_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na535_1_i) );
// C_AND////D      x51y46     80'h00_FE18_00_0000_0888_53FC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a536_1 ( .OUT(na536_1), .IN1(1'b1), .IN2(na88_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na88_1), .IN7(~na87_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a536_5 ( .OUT(na536_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na536_1) );
// C_MX2b/D///      x52y48     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a537_1 ( .OUT(na537_1_i), .IN1(1'b1), .IN2(~na536_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3717_2), .IN8(na538_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a537_2 ( .OUT(na537_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na537_1_i) );
// C_MX2b/D///      x48y40     80'h00_FE00_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a538_1 ( .OUT(na538_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4227_2), .IN5(1'b0), .IN6(na539_1), .IN7(1'b0), .IN8(na3716_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a538_2 ( .OUT(na538_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na538_1_i) );
// C_MX2b/D///      x45y38     80'h00_FE00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a539_1 ( .OUT(na539_1_i), .IN1(1'b1), .IN2(na536_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na540_1), .IN8(na3715_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a539_2 ( .OUT(na539_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na539_1_i) );
// C_MX2b/D///      x46y39     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a540_1 ( .OUT(na540_1_i), .IN1(1'b1), .IN2(~na536_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3714_1), .IN8(na541_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a540_2 ( .OUT(na540_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na540_1_i) );
// C_MX2b/D///      x46y40     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a541_1 ( .OUT(na541_1_i), .IN1(1'b1), .IN2(~na536_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3713_2), .IN8(na542_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a541_2 ( .OUT(na541_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na541_1_i) );
// C_MX2b/D///      x42y40     80'h00_FE00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a542_1 ( .OUT(na542_1_i), .IN1(1'b1), .IN2(na536_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na695_1), .IN8(na3712_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a542_2 ( .OUT(na542_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na542_1_i) );
// C_ORAND*/D//ORAND*/D      x61y51     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a543_1 ( .OUT(na543_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na543_2), .IN6(~na91_1), .IN7(~na2118_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a543_2 ( .OUT(na543_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na543_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a543_4 ( .OUT(na543_2_i), .IN1(~na545_1), .IN2(~na91_1), .IN3(~na2118_1), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a543_5 ( .OUT(na543_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na543_2_i) );
// C_ORAND*/D//ORAND*/D      x63y53     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a545_1 ( .OUT(na545_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na545_2), .IN6(~na91_1), .IN7(~na2120_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a545_2 ( .OUT(na545_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na545_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a545_4 ( .OUT(na545_2_i), .IN1(~na4231_2), .IN2(~na91_1), .IN3(~na2120_1), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a545_5 ( .OUT(na545_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na545_2_i) );
// C_ORAND*/D//ORAND*/D      x68y53     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a547_1 ( .OUT(na547_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4232_2), .IN6(~na91_1), .IN7(~na4501_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a547_2 ( .OUT(na547_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na547_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a547_4 ( .OUT(na547_2_i), .IN1(~na4233_2), .IN2(~na91_1), .IN3(~na4500_2), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a547_5 ( .OUT(na547_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na547_2_i) );
// C_ORAND*/D//ORAND*/D      x66y51     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a549_1 ( .OUT(na549_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4234_2), .IN6(~na91_1), .IN7(~na2124_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a549_2 ( .OUT(na549_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na549_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a549_4 ( .OUT(na549_2_i), .IN1(~na4235_2), .IN2(~na91_1), .IN3(~na2124_1), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a549_5 ( .OUT(na549_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na549_2_i) );
// C_ORAND*/D//ORAND*/D      x66y53     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a551_1 ( .OUT(na551_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4236_2), .IN6(~na91_1), .IN7(~na4482_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a551_2 ( .OUT(na551_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na551_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a551_4 ( .OUT(na551_2_i), .IN1(~na4237_2), .IN2(~na91_1), .IN3(~na4481_2), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a551_5 ( .OUT(na551_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na551_2_i) );
// C_ORAND*/D//ORAND*/D      x67y50     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a553_1 ( .OUT(na553_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4238_2), .IN6(~na91_1), .IN7(~na1889_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a553_2 ( .OUT(na553_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na553_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a553_4 ( .OUT(na553_2_i), .IN1(~na555_1), .IN2(~na91_1), .IN3(~na1889_1), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a553_5 ( .OUT(na553_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na553_2_i) );
// C_ORAND*/D//ORAND*/D      x67y51     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a555_1 ( .OUT(na555_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na555_2), .IN6(~na91_1), .IN7(~na1891_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a555_2 ( .OUT(na555_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na555_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a555_4 ( .OUT(na555_2_i), .IN1(~na557_1), .IN2(~na91_1), .IN3(~na1891_1), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a555_5 ( .OUT(na555_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na555_2_i) );
// C_ORAND*/D//ORAND*/D      x69y51     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a557_1 ( .OUT(na557_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na557_2), .IN6(~na91_1), .IN7(~na1893_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a557_2 ( .OUT(na557_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na557_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a557_4 ( .OUT(na557_2_i), .IN1(~na4243_2), .IN2(~na91_1), .IN3(~na1893_1), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a557_5 ( .OUT(na557_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na557_2_i) );
// C_ORAND*/D//ORAND*/D      x71y52     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a559_1 ( .OUT(na559_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4244_2), .IN6(~na91_1), .IN7(~na1862_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a559_2 ( .OUT(na559_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na559_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a559_4 ( .OUT(na559_2_i), .IN1(~na4245_2), .IN2(~na91_1), .IN3(~na1862_1), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a559_5 ( .OUT(na559_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na559_2_i) );
// C_ORAND*/D//ORAND*/D      x70y47     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a561_1 ( .OUT(na561_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4246_2), .IN6(~na91_1), .IN7(~na1864_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a561_2 ( .OUT(na561_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na561_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a561_4 ( .OUT(na561_2_i), .IN1(~na563_1), .IN2(~na91_1), .IN3(~na1864_1), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a561_5 ( .OUT(na561_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na561_2_i) );
// C_ORAND*/D//ORAND*/D      x67y49     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a563_1 ( .OUT(na563_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na563_2), .IN6(~na91_1), .IN7(~na1866_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a563_2 ( .OUT(na563_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na563_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a563_4 ( .OUT(na563_2_i), .IN1(~na565_1), .IN2(~na91_1), .IN3(~na1866_1), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a563_5 ( .OUT(na563_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na563_2_i) );
// C_ORAND*/D//ORAND*/D      x67y43     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a565_1 ( .OUT(na565_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na565_2), .IN6(~na91_1), .IN7(~na1868_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a565_2 ( .OUT(na565_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na565_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a565_4 ( .OUT(na565_2_i), .IN1(~na567_1), .IN2(~na91_1), .IN3(~na1868_1), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a565_5 ( .OUT(na565_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na565_2_i) );
// C_ORAND*/D//ORAND*/D      x63y43     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a567_1 ( .OUT(na567_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na567_2), .IN6(~na91_1), .IN7(~na3718_1),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a567_2 ( .OUT(na567_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na567_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a567_4 ( .OUT(na567_2_i), .IN1(~na569_1), .IN2(~na91_1), .IN3(~na3717_2), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a567_5 ( .OUT(na567_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na567_2_i) );
// C_ORAND*/D//ORAND*/D      x59y43     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a569_1 ( .OUT(na569_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na569_2), .IN6(~na91_1), .IN7(~na4617_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a569_2 ( .OUT(na569_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na569_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a569_4 ( .OUT(na569_2_i), .IN1(~na571_1), .IN2(~na91_1), .IN3(~na4616_2), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a569_5 ( .OUT(na569_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na569_2_i) );
// C_ORAND*/D//ORAND*/D      x59y45     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a571_1 ( .OUT(na571_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na571_2), .IN6(~na91_1), .IN7(~na3714_1),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a571_2 ( .OUT(na571_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na571_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a571_4 ( .OUT(na571_2_i), .IN1(~na573_1), .IN2(~na91_1), .IN3(~na3713_2), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a571_5 ( .OUT(na571_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na571_2_i) );
// C_ORAND*/D//ORAND*/D      x61y45     80'h00_F600_80_0000_0387_777B
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a573_1 ( .OUT(na573_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na573_2), .IN6(~na91_1), .IN7(~na4615_2),
                     .IN8(~na92_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a573_2 ( .OUT(na573_1), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na573_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a573_4 ( .OUT(na573_2_i), .IN1(na516_1), .IN2(~na91_1), .IN3(~na4614_2), .IN4(~na92_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a573_5 ( .OUT(na573_2), .CLK(na1739_1), .EN(~na1406_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na573_2_i) );
// C_ORAND////      x70y69     80'h00_0018_00_0000_0C88_E3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a575_1 ( .OUT(na575_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1986_1), .IN7(na38_1), .IN8(na3415_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/D      x48y55     80'h00_FE00_80_0000_0C0E_FFD0
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a576_4 ( .OUT(na576_2_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na3343_1), .IN4(na577_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a576_5 ( .OUT(na576_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na576_2_i) );
// C_AND////      x58y62     80'h00_0018_00_0000_0888_3C23
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a577_1 ( .OUT(na577_1), .IN1(1'b1), .IN2(~na1451_1), .IN3(na1991_1), .IN4(~na55_1), .IN5(1'b1), .IN6(na3196_1), .IN7(1'b1),
                     .IN8(~na55_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x52y57     80'h00_FE00_00_0040_0AA2_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a578_1 ( .OUT(na578_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na526_1), .IN5(1'b0), .IN6(~na428_1), .IN7(1'b0), .IN8(na1544_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a578_2 ( .OUT(na578_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na578_1_i) );
// C_MX2b/D///      x52y54     80'h00_FE00_00_0040_0AA2_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a579_1 ( .OUT(na579_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na526_1), .IN5(1'b0), .IN6(~na4096_2), .IN7(1'b0), .IN8(na1544_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a579_2 ( .OUT(na579_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na579_1_i) );
// C_ORAND/D///      x47y52     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a580_1 ( .OUT(na580_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4494_2), .IN6(~na3418_1), .IN7(~na3419_1),
                     .IN8(~na526_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a580_2 ( .OUT(na580_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na580_1_i) );
// C_///ORAND/D      x48y49     80'h00_FE00_80_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a582_4 ( .OUT(na582_2_i), .IN1(~na4495_2), .IN2(~na3418_1), .IN3(~na3422_1), .IN4(~na526_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a582_5 ( .OUT(na582_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na582_2_i) );
// C_ORAND/D///      x44y49     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a584_1 ( .OUT(na584_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2001_1), .IN6(~na3418_1), .IN7(~na3425_1),
                     .IN8(~na526_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a584_2 ( .OUT(na584_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na584_1_i) );
// C_ORAND/D///      x46y51     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a586_1 ( .OUT(na586_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4496_2), .IN6(~na3418_1), .IN7(~na3428_1),
                     .IN8(~na526_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a586_2 ( .OUT(na586_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na586_1_i) );
// C_ORAND/D///      x45y49     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a588_1 ( .OUT(na588_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2001_2), .IN6(~na3418_1), .IN7(~na3431_1),
                     .IN8(~na526_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a588_2 ( .OUT(na588_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na588_1_i) );
// C_MX2b/D///      x57y48     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a590_1 ( .OUT(na590_1_i), .IN1(1'b1), .IN2(na4223_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3432_1), .IN6(na3165_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a590_2 ( .OUT(na590_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na590_1_i) );
// C_MX2b/D///      x58y45     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a591_1 ( .OUT(na591_1_i), .IN1(1'b1), .IN2(na4223_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3433_2), .IN6(na3166_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a591_2 ( .OUT(na591_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na591_1_i) );
// C_MX2b/D///      x57y49     80'h00_FE00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a592_1 ( .OUT(na592_1_i), .IN1(1'b1), .IN2(~na4223_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3167_1), .IN6(na3434_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a592_2 ( .OUT(na592_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na592_1_i) );
// C_MX2b/D///      x55y45     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a593_1 ( .OUT(na593_1_i), .IN1(1'b1), .IN2(na4223_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3435_2), .IN6(na3168_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a593_2 ( .OUT(na593_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na593_1_i) );
// C_MX2b/D///      x56y54     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a594_1 ( .OUT(na594_1_i), .IN1(1'b1), .IN2(~na4223_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3169_1), .IN8(na3436_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a594_2 ( .OUT(na594_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na594_1_i) );
// C_MX2b/D///      x58y47     80'h00_FE00_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a595_1 ( .OUT(na595_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na526_1), .IN5(1'b0), .IN6(na3437_1), .IN7(1'b0), .IN8(na3170_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a595_2 ( .OUT(na595_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na595_1_i) );
// C_MX2b/D///      x54y50     80'h00_FE00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a596_1 ( .OUT(na596_1_i), .IN1(1'b1), .IN2(na4223_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3438_1), .IN8(na3171_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a596_2 ( .OUT(na596_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na596_1_i) );
// C_ORAND*////D      x66y68     80'h00_FE18_00_0000_0788_D55D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a597_1 ( .OUT(na597_1), .IN1(~na95_1), .IN2(na3440_1), .IN3(~na603_1), .IN4(1'b0), .IN5(~na95_2), .IN6(1'b0), .IN7(~na603_2),
                     .IN8(na614_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a597_5 ( .OUT(na597_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na597_1) );
// C_AND///AND/      x70y71     80'h00_0078_00_0000_0C88_12C3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a598_1 ( .OUT(na598_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3441_2), .IN6(~na1986_1), .IN7(~na4485_2),
                     .IN8(~na1985_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a598_4 ( .OUT(na598_2), .IN1(1'b1), .IN2(~na1986_1), .IN3(1'b1), .IN4(na1985_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x67y70     80'h00_0060_00_0000_0C06_FFB3
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a599_4 ( .OUT(na599_2), .IN1(1'b1), .IN2(na512_1), .IN3(~na3348_1), .IN4(na600_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x64y62     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a600_4 ( .OUT(na600_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1991_1), .IN4(na1984_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x64y73     80'h00_0078_00_0000_0C88_8C31
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a603_1 ( .OUT(na603_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3445_2), .IN7(na3451_2), .IN8(na56_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a603_4 ( .OUT(na603_2), .IN1(~na4489_2), .IN2(~na1993_2), .IN3(1'b1), .IN4(~na1990_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x66y78     80'h00_0018_00_0000_0C88_CBFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a605_1 ( .OUT(na605_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3447_2), .IN6(~na606_1), .IN7(1'b0), .IN8(na46_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x67y76     80'h00_0018_00_0040_0C68_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a606_1 ( .OUT(na606_1), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(na1990_1), .IN5(1'b1), .IN6(~na1989_2), .IN7(1'b1), .IN8(~na1990_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x67y77     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a607_1 ( .OUT(na607_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3448_1), .IN6(1'b0), .IN7(na3451_2), .IN8(~na2011_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x64y84     80'h00_0018_00_0000_0C66_6A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a612_1 ( .OUT(na612_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4080_2), .IN6(1'b0), .IN7(na613_2), .IN8(na1440_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x62y81     80'h00_0060_00_0000_0C08_FFA4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a613_4 ( .OUT(na613_2), .IN1(~na360_2), .IN2(na523_1), .IN3(na4086_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x68y66     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a614_1 ( .OUT(na614_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na575_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na3452_2), .IN7(1'b0), .IN8(~na1581_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x68y77     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a618_1 ( .OUT(na618_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1986_2), .IN7(1'b0), .IN8(na79_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x67y67     80'h00_0018_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a619_1 ( .OUT(na619_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4484_2), .IN5(na3164_1), .IN6(1'b0), .IN7(na3163_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x55y48     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a620_1 ( .OUT(na620_1_i), .IN1(1'b1), .IN2(na4223_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3458_2), .IN6(na3172_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a620_2 ( .OUT(na620_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na620_1_i) );
// C_MX2b////      x56y44     80'h00_0018_00_0040_0AA2_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a621_1 ( .OUT(na621_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na526_1), .IN5(1'b0), .IN6(~na89_2), .IN7(1'b0), .IN8(na1544_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x57y43     80'h00_0018_00_0040_0AA2_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a622_1 ( .OUT(na622_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na526_1), .IN5(1'b0), .IN6(~na89_1), .IN7(1'b0), .IN8(na1544_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x53y55     80'h00_0060_00_0000_0C08_FF75
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a623_4 ( .OUT(na623_2), .IN1(~na624_1), .IN2(1'b0), .IN3(~na3419_1), .IN4(~na526_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y55     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a624_1 ( .OUT(na624_1), .IN1(1'b1), .IN2(na536_1), .IN3(1'b1), .IN4(na526_1), .IN5(na496_1), .IN6(na1994_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x52y49     80'h00_0060_00_0000_0C08_FF73
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a625_4 ( .OUT(na625_2), .IN1(1'b0), .IN2(~na626_1), .IN3(~na3422_1), .IN4(~na526_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y56     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a626_1 ( .OUT(na626_1), .IN1(1'b1), .IN2(na536_1), .IN3(1'b1), .IN4(na526_1), .IN5(na499_1), .IN6(na1995_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x50y49     80'h00_0018_00_0000_0C88_75FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a627_1 ( .OUT(na627_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na628_1), .IN6(1'b0), .IN7(~na3425_1), .IN8(~na526_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y53     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a628_1 ( .OUT(na628_1), .IN1(1'b1), .IN2(na536_1), .IN3(1'b1), .IN4(na526_1), .IN5(na501_1), .IN6(na1996_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x48y51     80'h00_0018_00_0000_0C88_75FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a629_1 ( .OUT(na629_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na630_1), .IN6(1'b0), .IN7(~na3428_1), .IN8(~na526_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y51     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a630_1 ( .OUT(na630_1), .IN1(1'b1), .IN2(na536_1), .IN3(1'b1), .IN4(na526_1), .IN5(na503_1), .IN6(na1997_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x47y50     80'h00_0060_00_0000_0C08_FF75
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a631_4 ( .OUT(na631_2), .IN1(~na632_1), .IN2(1'b0), .IN3(~na3431_1), .IN4(~na526_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y47     80'h00_0018_00_0040_0A30_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a632_1 ( .OUT(na632_1), .IN1(1'b1), .IN2(na536_1), .IN3(1'b1), .IN4(na526_1), .IN5(na505_1), .IN6(na1998_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x17y78     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a633_1 ( .OUT(na633_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na634_1), .IN6(na633_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a633_2 ( .OUT(na633_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na633_1_i) );
// C_MX4b/D///      x19y75     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a634_1 ( .OUT(na634_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na634_1), .IN6(na635_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a634_2 ( .OUT(na634_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na634_1_i) );
// C_MX4b/D///      x19y76     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a635_1 ( .OUT(na635_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na1319_1), .IN6(na635_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a635_2 ( .OUT(na635_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na635_1_i) );
// C_ORAND////      x54y43     80'h00_0018_00_0000_0888_F5EA
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a636_1 ( .OUT(na636_1), .IN1(na3459_1), .IN2(1'b0), .IN3(na276_1), .IN4(na3462_1), .IN5(~na1473_2), .IN6(1'b0), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x51y55     80'h00_FE00_80_0000_0C08_FF2A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a638_4 ( .OUT(na638_2_i), .IN1(na1387_1), .IN2(1'b1), .IN3(na283_1), .IN4(~na282_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a638_5 ( .OUT(na638_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na638_2_i) );
// C_OR////D      x39y39     80'h00_FE18_00_0000_0EEE_50A0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a639_1 ( .OUT(na639_1), .IN1(1'b0), .IN2(1'b0), .IN3(na3463_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na636_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a639_5 ( .OUT(na639_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na639_1) );
// C_MX4b/D///      x19y78     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a640_1 ( .OUT(na640_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na641_1), .IN6(na640_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a640_2 ( .OUT(na640_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na640_1_i) );
// C_MX4b/D///      x21y77     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a641_1 ( .OUT(na641_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na641_1), .IN6(na642_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a641_2 ( .OUT(na641_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na641_1_i) );
// C_MX4b/D///      x23y78     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a642_1 ( .OUT(na642_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na674_1), .IN6(na642_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a642_2 ( .OUT(na642_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na642_1_i) );
// C_///AND/      x19y71     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a643_4 ( .OUT(na643_2), .IN1(1'b1), .IN2(~na405_2), .IN3(na317_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x16y69     80'h00_0018_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a644_1 ( .OUT(na644_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2_2), .IN7(~na318_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x36y70     80'h00_FE00_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a645_1 ( .OUT(na645_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3465_1), .IN6(~na3464_1), .IN7(~na1149_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a645_2 ( .OUT(na645_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na645_1_i) );
// C_MX4b/D///      x19y77     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a647_1 ( .OUT(na647_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na647_1), .IN6(na685_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a647_2 ( .OUT(na647_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na647_1_i) );
// C_MX2b/D///      x56y56     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a648_1 ( .OUT(na648_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na2358_1), .IN7(1'b0), .IN8(na649_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a648_2 ( .OUT(na648_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na648_1_i) );
// C_MX2b/D///      x56y52     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a649_1 ( .OUT(na649_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1741_2), .IN7(1'b0), .IN8(na650_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a649_2 ( .OUT(na649_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na649_1_i) );
// C_MX2b/D///      x56y50     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a650_1 ( .OUT(na650_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1741_1), .IN7(1'b0), .IN8(na651_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a650_2 ( .OUT(na650_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na650_1_i) );
// C_MX2b/D///      x60y48     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a651_1 ( .OUT(na651_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1743_2), .IN7(1'b0), .IN8(na652_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a651_2 ( .OUT(na651_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na651_1_i) );
// C_MX2b/D///      x56y46     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a652_1 ( .OUT(na652_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1743_1), .IN7(1'b0), .IN8(na658_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a652_2 ( .OUT(na652_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na652_1_i) );
// C_MX2b/D///      x56y55     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a653_1 ( .OUT(na653_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1882_2), .IN7(1'b0), .IN8(na654_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a653_2 ( .OUT(na653_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na653_1_i) );
// C_MX2b/D///      x54y52     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a654_1 ( .OUT(na654_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1882_1), .IN7(1'b0), .IN8(na655_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a654_2 ( .OUT(na654_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na654_1_i) );
// C_MX2b/D///      x58y48     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a655_1 ( .OUT(na655_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1884_2), .IN7(1'b0), .IN8(na656_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a655_2 ( .OUT(na655_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na655_1_i) );
// C_MX2b/D///      x58y46     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a656_1 ( .OUT(na656_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1884_1), .IN7(1'b0), .IN8(na657_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a656_2 ( .OUT(na656_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na656_1_i) );
// C_MX2b/D///      x50y44     80'h00_F600_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a657_1 ( .OUT(na657_1_i), .IN1(na1465_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3726_1), .IN8(na658_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a657_2 ( .OUT(na657_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na657_1_i) );
// C_MX2b/D///      x50y42     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a658_1 ( .OUT(na658_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4432_2), .IN5(na659_1), .IN6(1'b0), .IN7(na3725_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a658_2 ( .OUT(na658_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na658_1_i) );
// C_MX2b/D///      x47y41     80'h00_F600_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a659_1 ( .OUT(na659_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4432_2), .IN5(1'b0), .IN6(na660_1), .IN7(1'b0), .IN8(na3724_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a659_2 ( .OUT(na659_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na659_1_i) );
// C_MX2a/D///      x49y40     80'h00_F600_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a660_1 ( .OUT(na660_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na661_1), .IN4(na3723_2), .IN5(~na1465_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a660_2 ( .OUT(na660_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na660_1_i) );
// C_MX2b/D///      x48y41     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a661_1 ( .OUT(na661_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4432_2), .IN5(na662_1), .IN6(1'b0), .IN7(na3722_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a661_2 ( .OUT(na661_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na661_1_i) );
// C_MX2a/D///      x47y43     80'h00_F600_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a662_1 ( .OUT(na662_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na3721_2), .IN4(na1585_1), .IN5(na1465_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a662_2 ( .OUT(na662_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na662_1_i) );
// C_MX2b/D///      x55y52     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a663_1 ( .OUT(na663_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na2358_1), .IN7(1'b0), .IN8(na2230_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a663_2 ( .OUT(na663_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na663_1_i) );
// C_MX2a/D///      x59y56     80'h00_F600_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a664_1 ( .OUT(na664_1_i), .IN1(na665_1), .IN2(na1882_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1465_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a664_2 ( .OUT(na664_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na664_1_i) );
// C_MX2b/D///      x59y53     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a665_1 ( .OUT(na665_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1745_2), .IN7(1'b0), .IN8(na666_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a665_2 ( .OUT(na665_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na665_1_i) );
// C_MX2b/D///      x62y52     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a666_1 ( .OUT(na666_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1745_1), .IN7(1'b0), .IN8(na667_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a666_2 ( .OUT(na666_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na666_1_i) );
// C_MX2b/D///      x58y50     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a667_1 ( .OUT(na667_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1747_2), .IN7(1'b0), .IN8(na668_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a667_2 ( .OUT(na667_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na667_1_i) );
// C_MX2b/D///      x58y54     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a668_1 ( .OUT(na668_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1747_1), .IN7(1'b0), .IN8(na669_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a668_2 ( .OUT(na668_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na668_1_i) );
// C_MX2a/D///      x56y48     80'h00_F600_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a669_1 ( .OUT(na669_1_i), .IN1(na670_1), .IN2(na1878_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1465_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a669_2 ( .OUT(na669_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na669_1_i) );
// C_MX2b/D///      x61y49     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a670_1 ( .OUT(na670_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1878_1), .IN7(1'b0), .IN8(na671_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a670_2 ( .OUT(na670_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na670_1_i) );
// C_MX2a/D///      x54y48     80'h00_F600_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a671_1 ( .OUT(na671_1_i), .IN1(na672_1), .IN2(na1880_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1465_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a671_2 ( .OUT(na671_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na671_1_i) );
// C_MX2b/D///      x59y51     80'h00_F600_00_0040_0AA8_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a672_1 ( .OUT(na672_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4432_2), .IN5(1'b0), .IN6(na1880_1), .IN7(1'b0), .IN8(~na673_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a672_2 ( .OUT(na672_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na672_1_i) );
// C_MX2b////      x54y58     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a673_1 ( .OUT(na673_1), .IN1(na2229_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na653_1), .IN8(~na2230_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x25y77     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a674_1 ( .OUT(na674_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na674_1), .IN6(na4256_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a674_2 ( .OUT(na674_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na674_1_i) );
// C_MX2b/D///      x65y41     80'h00_FE00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a675_1 ( .OUT(na675_1_i), .IN1(1'b1), .IN2(~na4258_2), .IN3(1'b0), .IN4(1'b0), .IN5(na678_1), .IN6(na676_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a675_2 ( .OUT(na675_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na675_1_i) );
// C_MX2a////      x63y42     80'h00_0018_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a676_1 ( .OUT(na676_1), .IN1(na675_1), .IN2(na1747_1), .IN3(1'b0), .IN4(1'b0), .IN5(na275_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x62y48     80'h00_0060_00_0000_0C08_FF88
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a677_4 ( .OUT(na677_2), .IN1(na2229_1), .IN2(na2228_2), .IN3(na2223_2), .IN4(na4432_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x67y41     80'h00_FE00_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a678_1 ( .OUT(na678_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na677_2), .IN5(na680_1), .IN6(1'b0), .IN7(na679_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a678_2 ( .OUT(na678_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na678_1_i) );
// C_MX2b////      x58y43     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a679_1 ( .OUT(na679_1), .IN1(na275_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na678_1), .IN6(na1878_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x65y43     80'h00_FE00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a680_1 ( .OUT(na680_1_i), .IN1(1'b1), .IN2(~na4258_2), .IN3(1'b0), .IN4(1'b0), .IN5(na682_1), .IN6(na681_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a680_2 ( .OUT(na680_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na680_1_i) );
// C_MX2b////      x59y46     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a681_1 ( .OUT(na681_1), .IN1(na275_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na680_1), .IN6(na1878_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x65y45     80'h00_FE00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a682_1 ( .OUT(na682_1_i), .IN1(1'b1), .IN2(~na4258_2), .IN3(1'b0), .IN4(1'b0), .IN5(na684_1), .IN6(na683_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a682_2 ( .OUT(na682_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na682_1_i) );
// C_MX2a////      x57y46     80'h00_0018_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a683_1 ( .OUT(na683_1), .IN1(na682_1), .IN2(na1880_2), .IN3(1'b0), .IN4(1'b0), .IN5(na275_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x59y47     80'h00_FE00_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a684_1 ( .OUT(na684_1_i), .IN1(na275_2), .IN2(1'b1), .IN3(1'b1), .IN4(na677_2), .IN5(na684_1), .IN6(na1880_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a684_2 ( .OUT(na684_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na684_1_i) );
// C_MX4b/D///      x21y80     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a685_1 ( .OUT(na685_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na686_1), .IN6(na685_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a685_2 ( .OUT(na685_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na685_1_i) );
// C_MX4b/D///      x23y81     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a686_1 ( .OUT(na686_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na686_1), .IN6(na1318_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a686_2 ( .OUT(na686_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na686_1_i) );
// C_///AND/      x23y70     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a687_4 ( .OUT(na687_2), .IN1(1'b1), .IN2(na405_2), .IN3(1'b1), .IN4(na688_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x20y72     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a688_1 ( .OUT(na688_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4072_2), .IN7(1'b1), .IN8(~na26_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x16y74     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a689_1 ( .OUT(na689_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2_2), .IN7(na319_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x29y70     80'h00_FE00_00_0000_0C88_5DFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a690_1 ( .OUT(na690_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3466_2), .IN6(na3467_2), .IN7(~na1149_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a690_2 ( .OUT(na690_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na690_1_i) );
// C_MX4b/D///      x21y87     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a692_1 ( .OUT(na692_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na692_1), .IN6(na4259_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a692_2 ( .OUT(na692_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na692_1_i) );
// C_MX4b/D///      x23y87     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a693_1 ( .OUT(na693_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na693_1), .IN6(na694_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a693_2 ( .OUT(na693_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na693_1_i) );
// C_MX4b/D///      x19y88     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a694_1 ( .OUT(na694_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na696_1), .IN6(na694_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a694_2 ( .OUT(na694_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na694_1_i) );
// C_AND/D///      x44y39     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a695_1 ( .OUT(na695_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na536_1), .IN7(1'b1), .IN8(na3711_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a695_2 ( .OUT(na695_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na695_1_i) );
// C_MX4b/D///      x19y87     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a696_1 ( .OUT(na696_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na697_1), .IN6(na4260_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a696_2 ( .OUT(na696_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na696_1_i) );
// C_MX4b/D///      x21y85     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a697_1 ( .OUT(na697_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na697_1), .IN6(na710_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a697_2 ( .OUT(na697_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na697_1_i) );
// C_MX2a/D///      x25y37     80'h00_FE00_00_0040_0C05_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a698_1 ( .OUT(na698_1_i), .IN1(na699_1), .IN2(1'b0), .IN3(na3531_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na203_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a698_2 ( .OUT(na698_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na698_1_i) );
// C_MX2a/D///      x25y35     80'h00_FE00_00_0040_0C0A_CF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a699_1 ( .OUT(na699_1_i), .IN1(1'b0), .IN2(na700_1), .IN3(1'b0), .IN4(na3530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na203_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a699_2 ( .OUT(na699_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na699_1_i) );
// C_MX2a/D///      x25y40     80'h00_FE00_00_0040_0C0A_CF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a700_1 ( .OUT(na700_1_i), .IN1(1'b0), .IN2(na701_1), .IN3(1'b0), .IN4(na3529_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na203_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a700_2 ( .OUT(na700_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na700_1_i) );
// C_MX2b/D///      x33y40     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a701_1 ( .OUT(na701_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na203_2), .IN5(na702_1), .IN6(1'b0), .IN7(na3528_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a701_2 ( .OUT(na701_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na701_1_i) );
// C_MX2a/D///      x35y39     80'h00_FE00_00_0040_0C05_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a702_1 ( .OUT(na702_1_i), .IN1(na703_1), .IN2(1'b0), .IN3(na3527_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na203_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a702_2 ( .OUT(na702_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na702_1_i) );
// C_MX2b/D///      x35y37     80'h00_FE00_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a703_1 ( .OUT(na703_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na203_2), .IN5(1'b0), .IN6(na205_2), .IN7(1'b0), .IN8(na3526_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a703_2 ( .OUT(na703_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na703_1_i) );
// C_ANDXOR////D      x69y53     80'h00_FA18_00_0000_0666_3FB3
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a704_1 ( .OUT(na704_1), .IN1(1'b1), .IN2(na705_1), .IN3(~na3470_1), .IN4(na720_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1460_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a704_5 ( .OUT(na704_2), .CLK(na1739_1), .EN(na1459_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na704_1) );
// C_AND////      x63y62     80'h00_0018_00_0000_0C88_31FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a705_1 ( .OUT(na705_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na706_1), .IN6(~na3276_1), .IN7(1'b1), .IN8(~na4508_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x63y63     80'h00_0018_00_0000_0888_F9AA
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a706_1 ( .OUT(na706_1), .IN1(~na2229_1), .IN2(1'b0), .IN3(~na4263_2), .IN4(1'b0), .IN5(na2229_2), .IN6(na4505_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x59y61     80'h00_0018_00_0000_0C88_A2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a707_1 ( .OUT(na707_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na329_1), .IN6(~na295_1), .IN7(na262_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x65y55     80'h00_0060_00_0000_0C08_FFCD
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a708_4 ( .OUT(na708_2), .IN1(~na2229_1), .IN2(na3471_2), .IN3(1'b0), .IN4(na720_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x55y59     80'h00_F600_00_0040_0C03_0400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a709_1 ( .OUT(na709_1_i), .IN1(na704_1), .IN2(na2248_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na333_1), .IN6(na341_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a709_2 ( .OUT(na709_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na709_1_i) );
// C_MX4b/D///      x25y86     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a710_1 ( .OUT(na710_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na711_1), .IN6(na710_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a710_2 ( .OUT(na710_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na710_1_i) );
// C_MX4b/D///      x23y83     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a711_1 ( .OUT(na711_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na711_1), .IN6(na4264_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a711_2 ( .OUT(na711_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na711_1_i) );
// C_MX4b/D///      x25y83     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a712_1 ( .OUT(na712_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na712_1), .IN6(na1317_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a712_2 ( .OUT(na712_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na712_1_i) );
// C_ANDXOR/D//AND/D      x52y59     80'h00_FA00_80_0000_0C68_ECAF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a713_1 ( .OUT(na713_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na4175_2), .IN7(~na2223_2), .IN8(~na3472_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a713_2 ( .OUT(na713_1), .CLK(na1739_1), .EN(na1457_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na713_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a713_4 ( .OUT(na713_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na713_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a713_5 ( .OUT(na713_2), .CLK(na1739_1), .EN(na1457_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na713_2_i) );
// C_MX2b/D///      x48y38     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a714_1 ( .OUT(na714_1_i), .IN1(1'b1), .IN2(~na273_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3725_2), .IN8(na715_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a714_2 ( .OUT(na714_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na714_1_i) );
// C_MX2a/D///      x50y36     80'h00_FE00_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a715_1 ( .OUT(na715_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na716_1), .IN4(na3724_1), .IN5(1'b1), .IN6(na273_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a715_2 ( .OUT(na715_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na715_1_i) );
// C_MX2b/D///      x46y35     80'h00_FE00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a716_1 ( .OUT(na716_1_i), .IN1(1'b1), .IN2(na273_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na717_1), .IN8(na3723_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a716_2 ( .OUT(na716_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na716_1_i) );
// C_MX2a/D///      x46y37     80'h00_FE00_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a717_1 ( .OUT(na717_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na3722_1), .IN4(na718_1), .IN5(1'b1), .IN6(~na273_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a717_2 ( .OUT(na717_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na717_1_i) );
// C_MX2b/D///      x46y38     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a718_1 ( .OUT(na718_1_i), .IN1(1'b1), .IN2(~na273_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3721_2), .IN8(na719_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a718_2 ( .OUT(na718_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na718_1_i) );
// C_MX2a/D///      x44y38     80'h00_FE00_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a719_1 ( .OUT(na719_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na269_2), .IN4(na3720_1), .IN5(1'b1), .IN6(na273_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a719_2 ( .OUT(na719_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na719_1_i) );
// C_MX2b/D///      x60y50     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a720_1 ( .OUT(na720_1_i), .IN1(1'b1), .IN2(~na273_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3726_1), .IN8(na721_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a720_2 ( .OUT(na720_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na720_1_i) );
// C_MX2b/D///      x50y38     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a721_1 ( .OUT(na721_1_i), .IN1(1'b1), .IN2(~na273_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3725_2), .IN8(na722_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a721_2 ( .OUT(na721_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na721_1_i) );
// C_MX2a/D///      x52y36     80'h00_FE00_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a722_1 ( .OUT(na722_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na723_1), .IN4(na3724_1), .IN5(1'b1), .IN6(na273_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a722_2 ( .OUT(na722_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na722_1_i) );
// C_MX2b/D///      x48y37     80'h00_FE00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a723_1 ( .OUT(na723_1_i), .IN1(1'b1), .IN2(na273_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na724_1), .IN8(na3723_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a723_2 ( .OUT(na723_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na723_1_i) );
// C_MX2a/D///      x42y39     80'h00_FE00_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a724_1 ( .OUT(na724_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na3722_1), .IN4(na725_1), .IN5(1'b1), .IN6(~na273_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a724_2 ( .OUT(na724_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na724_1_i) );
// C_MX2b/D///      x42y38     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a725_1 ( .OUT(na725_1_i), .IN1(1'b1), .IN2(~na273_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3721_2), .IN8(na726_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a725_2 ( .OUT(na725_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na725_1_i) );
// C_MX2b/D///      x44y36     80'h00_FE00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a726_1 ( .OUT(na726_1_i), .IN1(1'b1), .IN2(na273_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na272_1), .IN8(na3720_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a726_2 ( .OUT(na726_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na726_1_i) );
// C_MX4b/D///      x19y85     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a727_1 ( .OUT(na727_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na760_1), .IN6(na4266_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a727_2 ( .OUT(na727_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na727_1_i) );
// C_ORAND*/D//ORAND*/D      x64y42     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a728_1 ( .OUT(na728_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na2352_2), .IN7(~na4268_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a728_2 ( .OUT(na728_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na728_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a728_4 ( .OUT(na728_2_i), .IN1(~na337_2), .IN2(~na2352_1), .IN3(~na730_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a728_5 ( .OUT(na728_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na728_2_i) );
// C_ORAND*/D//ORAND*/D      x62y41     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a730_1 ( .OUT(na730_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na2354_2), .IN7(~na730_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a730_2 ( .OUT(na730_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na730_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a730_4 ( .OUT(na730_2_i), .IN1(~na337_2), .IN2(~na2354_1), .IN3(~na732_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a730_5 ( .OUT(na730_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na730_2_i) );
// C_ORAND*/D//ORAND*/D      x62y43     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a732_1 ( .OUT(na732_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na2356_2), .IN7(~na732_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a732_2 ( .OUT(na732_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na732_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a732_4 ( .OUT(na732_2_i), .IN1(~na337_2), .IN2(~na2356_1), .IN3(~na4269_2), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a732_5 ( .OUT(na732_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na732_2_i) );
// C_ORAND*/D//ORAND*/D      x61y43     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a734_1 ( .OUT(na734_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na2358_2), .IN7(~na4270_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a734_2 ( .OUT(na734_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na734_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a734_4 ( .OUT(na734_2_i), .IN1(~na337_2), .IN2(~na2358_1), .IN3(~na736_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a734_5 ( .OUT(na734_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na734_2_i) );
// C_ORAND*/D//ORAND*/D      x66y41     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a736_1 ( .OUT(na736_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na1741_2), .IN7(~na736_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a736_2 ( .OUT(na736_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na736_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a736_4 ( .OUT(na736_2_i), .IN1(~na337_2), .IN2(~na1741_1), .IN3(~na738_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a736_5 ( .OUT(na736_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na736_2_i) );
// C_ORAND*/D//ORAND*/D      x68y39     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a738_1 ( .OUT(na738_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na1743_2), .IN7(~na738_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a738_2 ( .OUT(na738_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na738_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a738_4 ( .OUT(na738_2_i), .IN1(~na337_2), .IN2(~na1743_1), .IN3(~na740_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a738_5 ( .OUT(na738_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na738_2_i) );
// C_ORAND*/D//ORAND*/D      x72y39     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a740_1 ( .OUT(na740_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na1745_2), .IN7(~na740_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a740_2 ( .OUT(na740_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na740_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a740_4 ( .OUT(na740_2_i), .IN1(~na337_2), .IN2(~na1745_1), .IN3(~na742_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a740_5 ( .OUT(na740_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na740_2_i) );
// C_ORAND*/D//ORAND*/D      x70y41     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a742_1 ( .OUT(na742_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na1747_2), .IN7(~na742_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a742_2 ( .OUT(na742_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na742_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a742_4 ( .OUT(na742_2_i), .IN1(~na337_2), .IN2(~na1747_1), .IN3(~na744_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a742_5 ( .OUT(na742_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na742_2_i) );
// C_ORAND*/D//ORAND*/D      x70y37     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a744_1 ( .OUT(na744_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na1878_2), .IN7(~na744_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a744_2 ( .OUT(na744_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na744_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a744_4 ( .OUT(na744_2_i), .IN1(~na337_2), .IN2(~na1878_1), .IN3(~na746_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a744_5 ( .OUT(na744_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na744_2_i) );
// C_ORAND*/D//ORAND*/D      x68y37     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a746_1 ( .OUT(na746_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na1880_2), .IN7(~na746_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a746_2 ( .OUT(na746_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na746_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a746_4 ( .OUT(na746_2_i), .IN1(~na337_2), .IN2(~na1880_1), .IN3(~na748_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a746_5 ( .OUT(na746_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na746_2_i) );
// C_ORAND*/D//ORAND*/D      x70y39     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a748_1 ( .OUT(na748_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na1882_2), .IN7(~na748_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a748_2 ( .OUT(na748_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na748_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a748_4 ( .OUT(na748_2_i), .IN1(~na337_2), .IN2(~na1882_1), .IN3(~na750_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a748_5 ( .OUT(na748_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na748_2_i) );
// C_ORAND*/D//ORAND*/D      x66y39     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a750_1 ( .OUT(na750_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na1884_2), .IN7(~na750_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a750_2 ( .OUT(na750_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na750_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a750_4 ( .OUT(na750_2_i), .IN1(~na337_2), .IN2(~na1884_1), .IN3(~na4283_2), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a750_5 ( .OUT(na750_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na750_2_i) );
// C_ORAND*/D//ORAND*/D      x65y35     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a752_1 ( .OUT(na752_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na4625_2), .IN7(~na4284_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a752_2 ( .OUT(na752_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na752_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a752_4 ( .OUT(na752_2_i), .IN1(~na337_2), .IN2(~na4624_2), .IN3(~na4285_2), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a752_5 ( .OUT(na752_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na752_2_i) );
// C_ORAND*/D//ORAND*/D      x59y38     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a754_1 ( .OUT(na754_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na4623_2), .IN7(~na4286_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a754_2 ( .OUT(na754_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na754_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a754_4 ( .OUT(na754_2_i), .IN1(~na337_2), .IN2(~na4622_2), .IN3(~na4287_2), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a754_5 ( .OUT(na754_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na754_2_i) );
// C_ORAND*/D//ORAND*/D      x61y38     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a756_1 ( .OUT(na756_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na4621_2), .IN7(~na4288_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a756_2 ( .OUT(na756_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na756_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a756_4 ( .OUT(na756_2_i), .IN1(~na337_2), .IN2(~na4620_2), .IN3(~na758_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a756_5 ( .OUT(na756_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na756_2_i) );
// C_ORAND*/D//ORAND*/D      x58y35     80'h00_F600_80_0000_0387_77B7
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a758_1 ( .OUT(na758_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na337_2), .IN6(~na4619_2), .IN7(~na758_2),
                     .IN8(~na336_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a758_2 ( .OUT(na758_1), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na758_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a758_4 ( .OUT(na758_2_i), .IN1(~na337_2), .IN2(~na4618_2), .IN3(na354_1), .IN4(~na336_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a758_5 ( .OUT(na758_2), .CLK(na1739_1), .EN(~na1407_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na758_2_i) );
// C_MX4b/D///      x23y85     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a760_1 ( .OUT(na760_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na760_1), .IN6(na4291_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a760_2 ( .OUT(na760_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na760_1_i) );
// C_///ORAND/      x67y53     80'h00_0060_00_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a761_4 ( .OUT(na761_2), .IN1(na4161_2), .IN2(na3539_1), .IN3(~na2223_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x21y81     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a762_1 ( .OUT(na762_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na762_1), .IN6(na814_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a762_2 ( .OUT(na762_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na762_1_i) );
// C_///OR/D      x43y47     80'h00_FE00_80_0000_0C0E_FFA5
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a763_4 ( .OUT(na763_2_i), .IN1(~na3459_1), .IN2(1'b0), .IN3(na764_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a763_5 ( .OUT(na763_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na763_2_i) );
// C_AND////      x58y51     80'h00_0018_00_0000_0888_4CF4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a764_1 ( .OUT(na764_1), .IN1(~na1473_2), .IN2(na2228_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3461_1), .IN7(~na276_1),
                     .IN8(na3162_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x50y46     80'h00_FE00_00_0040_0AA8_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a765_1 ( .OUT(na765_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na636_1), .IN4(1'b1), .IN5(1'b0), .IN6(na1542_2), .IN7(1'b0), .IN8(~na4418_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a765_2 ( .OUT(na765_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na765_1_i) );
// C_MX2b/D///      x50y45     80'h00_FE00_00_0040_0AA8_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a766_1 ( .OUT(na766_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na636_1), .IN4(1'b1), .IN5(1'b0), .IN6(na1542_1), .IN7(1'b0), .IN8(~na284_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a766_2 ( .OUT(na766_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na766_1_i) );
// C_ORAND/D///      x48y48     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a767_1 ( .OUT(na767_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3542_1), .IN6(~na4513_2), .IN7(~na636_1),
                     .IN8(~na3543_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a767_2 ( .OUT(na767_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na767_1_i) );
// C_ORAND/D///      x44y47     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a769_1 ( .OUT(na769_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3542_1), .IN6(~na4514_2), .IN7(~na636_1),
                     .IN8(~na3546_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a769_2 ( .OUT(na769_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na769_1_i) );
// C_///ORAND/D      x46y48     80'h00_FE00_80_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a771_4 ( .OUT(na771_2_i), .IN1(~na3542_1), .IN2(~na2238_1), .IN3(~na636_1), .IN4(~na3549_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a771_5 ( .OUT(na771_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na771_2_i) );
// C_///ORAND/D      x48y48     80'h00_FE00_80_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a773_4 ( .OUT(na773_2_i), .IN1(~na3542_1), .IN2(~na4515_2), .IN3(~na636_1), .IN4(~na3552_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a773_5 ( .OUT(na773_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na773_2_i) );
// C_///ORAND/D      x44y47     80'h00_FE00_80_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a775_4 ( .OUT(na775_2_i), .IN1(~na3542_1), .IN2(~na2238_2), .IN3(~na636_1), .IN4(~na3555_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a775_5 ( .OUT(na775_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na775_2_i) );
// C_MX2b/D///      x56y38     80'h00_FE00_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a777_1 ( .OUT(na777_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na636_1), .IN4(1'b1), .IN5(na3556_2), .IN6(1'b0), .IN7(na3177_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a777_2 ( .OUT(na777_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na777_1_i) );
// C_MX2b/D///      x56y35     80'h00_FE00_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a778_1 ( .OUT(na778_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na636_1), .IN4(1'b1), .IN5(1'b0), .IN6(na3557_2), .IN7(1'b0), .IN8(na3178_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a778_2 ( .OUT(na778_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na778_1_i) );
// C_MX2b/D///      x52y37     80'h00_FE00_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a779_1 ( .OUT(na779_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na636_1), .IN4(1'b1), .IN5(na3558_2), .IN6(1'b0), .IN7(na3179_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a779_2 ( .OUT(na779_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na779_1_i) );
// C_MX2b/D///      x55y37     80'h00_FE00_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a780_1 ( .OUT(na780_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na636_1), .IN4(1'b1), .IN5(1'b0), .IN6(na3559_1), .IN7(1'b0), .IN8(na3180_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a780_2 ( .OUT(na780_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na780_1_i) );
// C_MX2b/D///      x56y42     80'h00_FE00_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a781_1 ( .OUT(na781_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(~na636_1), .IN4(1'b1), .IN5(na3181_1), .IN6(1'b0), .IN7(na3560_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a781_2 ( .OUT(na781_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na781_1_i) );
// C_MX2b/D///      x56y39     80'h00_FE00_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a782_1 ( .OUT(na782_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(na636_1), .IN4(1'b1), .IN5(1'b0), .IN6(na3561_1), .IN7(1'b0), .IN8(na3182_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a782_2 ( .OUT(na782_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na782_1_i) );
// C_MX2b/D///      x52y39     80'h00_FE00_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a783_1 ( .OUT(na783_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na636_1), .IN4(1'b1), .IN5(na3562_2), .IN6(1'b0), .IN7(na3183_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a783_2 ( .OUT(na783_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na783_1_i) );
// C_ORAND*////D      x62y55     80'h00_FE18_00_0000_0788_D35B
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a784_1 ( .OUT(na784_1), .IN1(na3564_1), .IN2(~na341_1), .IN3(~na790_1), .IN4(1'b0), .IN5(1'b0), .IN6(~na341_2), .IN7(~na790_2),
                     .IN8(na792_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a784_5 ( .OUT(na784_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na784_1) );
// C_AND///AND/      x67y55     80'h00_0078_00_0000_0C88_145A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a785_1 ( .OUT(na785_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2222_1), .IN6(na3565_2), .IN7(~na2223_1),
                     .IN8(~na4504_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a785_4 ( .OUT(na785_2), .IN1(na2222_1), .IN2(1'b1), .IN3(~na2223_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x61y54     80'h00_0018_00_0000_0C66_5D00
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a786_1 ( .OUT(na786_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na787_1), .IN6(~na4604_2), .IN7(na353_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x59y49     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a787_1 ( .OUT(na787_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2228_1), .IN7(1'b1), .IN8(na2221_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x54y61     80'h00_0078_00_0000_0C88_8A31
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a790_1 ( .OUT(na790_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3278_2), .IN6(1'b1), .IN7(na326_1), .IN8(na3272_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a790_4 ( .OUT(na790_2), .IN1(~na2229_1), .IN2(~na2228_2), .IN3(1'b1), .IN4(~na4511_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y52     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a792_1 ( .OUT(na792_1), .IN1(~na761_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3570_2), .IN6(~na1587_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x57y58     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a796_4 ( .OUT(na796_2), .IN1(1'b0), .IN2(na268_2), .IN3(na2223_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x70y55     80'h00_0018_00_0040_0A50_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a797_1 ( .OUT(na797_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2223_1), .IN4(1'b1), .IN5(na3175_1), .IN6(1'b0), .IN7(na3176_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x53y39     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a798_1 ( .OUT(na798_1_i), .IN1(1'b1), .IN2(na4255_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3576_2), .IN6(na3184_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a798_2 ( .OUT(na798_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na798_1_i) );
// C_MX2b////      x59y36     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a799_1 ( .OUT(na799_1), .IN1(1'b1), .IN2(na4255_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na4150_2), .IN6(na1542_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x60y35     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a800_1 ( .OUT(na800_1), .IN1(1'b1), .IN2(na4255_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na4149_2), .IN6(na1542_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x49y43     80'h00_0060_00_0000_0C08_FF75
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a801_4 ( .OUT(na801_2), .IN1(~na802_1), .IN2(1'b0), .IN3(~na636_1), .IN4(~na3543_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y41     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a802_1 ( .OUT(na802_1), .IN1(1'b1), .IN2(na273_1), .IN3(na636_1), .IN4(1'b1), .IN5(na675_1), .IN6(na2231_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x50y43     80'h00_0018_00_0000_0C88_73FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a803_1 ( .OUT(na803_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na804_1), .IN7(~na636_1), .IN8(~na3546_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y44     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a804_1 ( .OUT(na804_1), .IN1(1'b1), .IN2(na273_1), .IN3(na636_1), .IN4(1'b1), .IN5(na678_1), .IN6(na2232_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x49y43     80'h00_0018_00_0000_0C88_75FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a805_1 ( .OUT(na805_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na806_1), .IN6(1'b0), .IN7(~na636_1), .IN8(~na3549_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y39     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a806_1 ( .OUT(na806_1), .IN1(1'b1), .IN2(na273_1), .IN3(na636_1), .IN4(1'b1), .IN5(na680_1), .IN6(na2233_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x48y43     80'h00_0060_00_0000_0C08_FF75
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a807_4 ( .OUT(na807_2), .IN1(~na808_1), .IN2(1'b0), .IN3(~na636_1), .IN4(~na3552_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y43     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a808_1 ( .OUT(na808_1), .IN1(1'b1), .IN2(na273_1), .IN3(na636_1), .IN4(1'b1), .IN5(na682_1), .IN6(na2234_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x48y43     80'h00_0018_00_0000_0C88_73FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a809_1 ( .OUT(na809_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na810_1), .IN7(~na636_1), .IN8(~na3555_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x51y40     80'h00_0018_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a810_1 ( .OUT(na810_1), .IN1(1'b1), .IN2(na273_1), .IN3(na636_1), .IN4(1'b1), .IN5(na684_1), .IN6(na2235_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x48y85     80'h00_FE00_00_0040_0AC8_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a811_1 ( .OUT(na811_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na811_1), .IN8(~na812_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a811_2 ( .OUT(na811_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na811_1_i) );
// C_MX2b////      x58y86     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a812_1 ( .OUT(na812_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1085_1), .IN5(1'b0), .IN6(~na813_1), .IN7(1'b0), .IN8(~na612_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x63y78     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a813_1 ( .OUT(na813_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3445_2), .IN7(1'b1), .IN8(na56_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x23y80     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a814_1 ( .OUT(na814_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na815_1), .IN6(na814_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a814_2 ( .OUT(na814_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na814_1_i) );
// C_MX4b/D///      x23y79     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a815_1 ( .OUT(na815_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na816_1), .IN6(na4292_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a815_2 ( .OUT(na815_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na815_1_i) );
// C_MX4b/D///      x25y81     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a816_1 ( .OUT(na816_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na816_1), .IN6(na4294_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a816_2 ( .OUT(na816_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na816_1_i) );
// C_ORAND////      x47y76     80'h00_0018_00_0000_0888_5FAD
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a817_1 ( .OUT(na817_1), .IN1(~na4610_2), .IN2(na219_2), .IN3(na4609_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(~na1517_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x45y84     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a819_4 ( .OUT(na819_2), .IN1(1'b1), .IN2(~na219_2), .IN3(na3580_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y83     80'h00_0018_00_0000_0888_53A1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a820_1 ( .OUT(na820_1), .IN1(~na2712_2), .IN2(~na232_1), .IN3(na1340_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na4553_2), .IN7(~na2713_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x51y85     80'h00_FE00_00_0000_0C88_2CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a821_1 ( .OUT(na821_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1325_1), .IN7(na1326_1), .IN8(~na409_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a821_2 ( .OUT(na821_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na821_1_i) );
// C_OR////D      x33y60     80'h00_FE18_00_0000_0EEE_C003
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a822_1 ( .OUT(na822_1), .IN1(1'b0), .IN2(~na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3582_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a822_5 ( .OUT(na822_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na822_1) );
// C_MX4b/D///      x28y82     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a823_1 ( .OUT(na823_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1309_1),
                     .IN8(na823_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a823_2 ( .OUT(na823_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na823_1_i) );
// C_AND/D///      x69y90     80'h00_FE00_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a825_1 ( .OUT(na825_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1633_1), .IN6(1'b1), .IN7(~na443_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a825_2 ( .OUT(na825_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na825_1_i) );
// C_AND/D//AND/D      x70y90     80'h00_FE00_80_0000_0C88_5A1F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a826_1 ( .OUT(na826_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1633_2), .IN6(1'b1), .IN7(~na443_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a826_2 ( .OUT(na826_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na826_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a826_4 ( .OUT(na826_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na443_1), .IN4(~na826_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a826_5 ( .OUT(na826_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na826_2_i) );
// C_MX2b/D///      x23y52     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a827_1 ( .OUT(na827_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na828_1), .IN6(1'b0), .IN7(na2599_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a827_2 ( .OUT(na827_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na827_1_i) );
// C_MX2b/D///      x23y49     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a828_1 ( .OUT(na828_1_i), .IN1(1'b1), .IN2(na1487_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1819_2), .IN8(na829_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a828_2 ( .OUT(na828_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na828_1_i) );
// C_MX2b/D///      x22y48     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a829_1 ( .OUT(na829_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na830_1), .IN6(1'b0), .IN7(na1819_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a829_2 ( .OUT(na829_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na829_1_i) );
// C_MX2b/D///      x21y47     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a830_1 ( .OUT(na830_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na831_1), .IN6(1'b0), .IN7(na1821_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a830_2 ( .OUT(na830_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na830_1_i) );
// C_MX2b/D///      x21y45     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a831_1 ( .OUT(na831_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na837_1), .IN6(1'b0), .IN7(na1821_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a831_2 ( .OUT(na831_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na831_1_i) );
// C_MX2b/D///      x21y53     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a832_1 ( .OUT(na832_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na833_1), .IN6(1'b0), .IN7(na1815_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a832_2 ( .OUT(na832_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na832_1_i) );
// C_MX2b/D///      x27y49     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a833_1 ( .OUT(na833_1_i), .IN1(1'b1), .IN2(na1487_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1815_1), .IN8(na834_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a833_2 ( .OUT(na833_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na833_1_i) );
// C_MX2b/D///      x24y52     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a834_1 ( .OUT(na834_1_i), .IN1(1'b1), .IN2(na1487_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1817_2), .IN8(na835_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a834_2 ( .OUT(na834_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na834_1_i) );
// C_MX2b/D///      x24y46     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a835_1 ( .OUT(na835_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na836_1), .IN6(1'b0), .IN7(na1817_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a835_2 ( .OUT(na835_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na835_1_i) );
// C_MX2b/D///      x21y41     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a836_1 ( .OUT(na836_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na837_1), .IN6(1'b0), .IN7(na3532_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a836_2 ( .OUT(na836_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na836_1_i) );
// C_MX2b/D///      x21y39     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a837_1 ( .OUT(na837_1_i), .IN1(1'b1), .IN2(na1487_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3531_2), .IN8(na838_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a837_2 ( .OUT(na837_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na837_1_i) );
// C_MX2b/D///      x24y40     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a838_1 ( .OUT(na838_1_i), .IN1(1'b1), .IN2(~na1487_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na839_1), .IN8(na3530_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a838_2 ( .OUT(na838_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na838_1_i) );
// C_MX2b/D///      x22y37     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a839_1 ( .OUT(na839_1_i), .IN1(1'b1), .IN2(~na1487_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na840_1), .IN8(na3529_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a839_2 ( .OUT(na839_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na839_1_i) );
// C_MX2b/D///      x24y37     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a840_1 ( .OUT(na840_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na841_1), .IN6(1'b0), .IN7(na3528_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a840_2 ( .OUT(na840_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na840_1_i) );
// C_MX2b/D///      x23y41     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a841_1 ( .OUT(na841_1_i), .IN1(1'b1), .IN2(na1487_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3527_2), .IN8(na1591_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a841_2 ( .OUT(na841_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na841_1_i) );
// C_MX2b/D///      x19y46     80'h00_F600_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a842_1 ( .OUT(na842_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4442_2), .IN5(na4543_2), .IN6(1'b0), .IN7(na2481_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a842_2 ( .OUT(na842_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na842_1_i) );
// C_MX2b/D///      x19y53     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a843_1 ( .OUT(na843_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na844_1), .IN6(1'b0), .IN7(na1815_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a843_2 ( .OUT(na843_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na843_1_i) );
// C_MX2b/D///      x25y57     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a844_1 ( .OUT(na844_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na845_1), .IN6(1'b0), .IN7(na1823_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a844_2 ( .OUT(na844_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na844_1_i) );
// C_MX2b/D///      x29y55     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a845_1 ( .OUT(na845_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na846_1), .IN6(1'b0), .IN7(na1823_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a845_2 ( .OUT(na845_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na845_1_i) );
// C_MX2b/D///      x23y53     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a846_1 ( .OUT(na846_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na847_1), .IN6(1'b0), .IN7(na1825_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a846_2 ( .OUT(na846_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na846_1_i) );
// C_MX2b/D///      x27y53     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a847_1 ( .OUT(na847_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na848_1), .IN6(1'b0), .IN7(na1825_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a847_2 ( .OUT(na847_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na847_1_i) );
// C_MX2b/D///      x27y51     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a848_1 ( .OUT(na848_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na849_1), .IN6(1'b0), .IN7(na1811_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a848_2 ( .OUT(na848_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na848_1_i) );
// C_MX2a/D///      x29y53     80'h00_F600_00_0040_0C05_3000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a849_1 ( .OUT(na849_1_i), .IN1(na850_1), .IN2(1'b0), .IN3(na1811_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na4442_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a849_2 ( .OUT(na849_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na849_1_i) );
// C_MX2b/D///      x27y55     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a850_1 ( .OUT(na850_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(na851_1), .IN6(1'b0), .IN7(na1813_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a850_2 ( .OUT(na850_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na850_1_i) );
// C_MX2b/D///      x23y47     80'h00_F600_00_0040_0A51_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a851_1 ( .OUT(na851_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4442_2), .IN5(~na852_1), .IN6(1'b0), .IN7(na1813_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a851_2 ( .OUT(na851_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na851_1_i) );
// C_MX2b////      x19y47     80'h00_0018_00_0040_0A55_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a852_1 ( .OUT(na852_1), .IN1(1'b0), .IN2(1'b0), .IN3(na2481_2), .IN4(1'b1), .IN5(~na832_1), .IN6(1'b0), .IN7(~na2481_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x28y56     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a853_1 ( .OUT(na853_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na855_1), .IN5(na854_1), .IN6(1'b0), .IN7(na856_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a853_2 ( .OUT(na853_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na853_1_i) );
// C_MX2a////      x29y51     80'h00_0018_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a854_1 ( .OUT(na854_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1825_1), .IN4(na853_1), .IN5(~na121_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x26y54     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a855_1 ( .OUT(na855_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4522_2), .IN6(na2478_1), .IN7(na2481_2), .IN8(na4442_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x30y55     80'h00_FE00_00_0040_0C05_3000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a856_1 ( .OUT(na856_1_i), .IN1(na858_1), .IN2(1'b0), .IN3(na857_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na855_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a856_2 ( .OUT(na856_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na856_1_i) );
// C_MX2b////      x30y51     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a857_1 ( .OUT(na857_1), .IN1(na121_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na856_1), .IN8(na4479_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x31y55     80'h00_FE00_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a858_1 ( .OUT(na858_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na855_1), .IN5(1'b0), .IN6(na859_1), .IN7(1'b0), .IN8(na860_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a858_2 ( .OUT(na858_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na858_1_i) );
// C_MX2a////      x27y50     80'h00_0018_00_0040_0C03_0A00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a859_1 ( .OUT(na859_1), .IN1(na858_1), .IN2(na4478_2), .IN3(1'b0), .IN4(1'b0), .IN5(na121_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x30y56     80'h00_FE00_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a860_1 ( .OUT(na860_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na855_1), .IN5(1'b0), .IN6(na861_1), .IN7(1'b0), .IN8(na862_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a860_2 ( .OUT(na860_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na860_1_i) );
// C_MX2a////      x29y50     80'h00_0018_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a861_1 ( .OUT(na861_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1813_2), .IN4(na860_1), .IN5(~na121_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x30y52     80'h00_FE00_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a862_1 ( .OUT(na862_1_i), .IN1(~na121_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na855_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1813_1),
                     .IN8(na862_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a862_2 ( .OUT(na862_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na862_1_i) );
// C_MX2b/D///      x26y52     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a864_1 ( .OUT(na864_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na203_1), .IN5(na865_1), .IN6(1'b0), .IN7(na3532_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a864_2 ( .OUT(na864_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na864_1_i) );
// C_MX2b/D///      x23y39     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a865_1 ( .OUT(na865_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na203_1), .IN5(na866_1), .IN6(1'b0), .IN7(na3531_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a865_2 ( .OUT(na865_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na865_1_i) );
// C_MX2b/D///      x23y37     80'h00_FE00_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a866_1 ( .OUT(na866_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na203_1), .IN5(1'b0), .IN6(na867_1), .IN7(1'b0), .IN8(na3530_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a866_2 ( .OUT(na866_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na866_1_i) );
// C_MX2a/D///      x23y36     80'h00_FE00_00_0040_0C0A_CF00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a867_1 ( .OUT(na867_1_i), .IN1(1'b0), .IN2(na868_1), .IN3(1'b0), .IN4(na3529_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na203_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a867_2 ( .OUT(na867_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na867_1_i) );
// C_MX2b/D///      x27y40     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a868_1 ( .OUT(na868_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na203_1), .IN5(na869_1), .IN6(1'b0), .IN7(na3528_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a868_2 ( .OUT(na868_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na868_1_i) );
// C_MX2a/D///      x27y37     80'h00_FE00_00_0040_0C05_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a869_1 ( .OUT(na869_1_i), .IN1(na870_1), .IN2(1'b0), .IN3(na3527_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na203_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a869_2 ( .OUT(na869_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na869_1_i) );
// C_MX2b/D///      x29y35     80'h00_FE00_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a870_1 ( .OUT(na870_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na203_1), .IN5(1'b0), .IN6(na202_1), .IN7(1'b0), .IN8(na3526_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a870_2 ( .OUT(na870_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na870_1_i) );
// C_MX2b/D///      x40y56     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a871_1 ( .OUT(na871_1_i), .IN1(~na399_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3423_2), .IN8(na872_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a871_2 ( .OUT(na871_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na871_1_i) );
// C_MX2b/D///      x40y52     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a872_1 ( .OUT(na872_1_i), .IN1(na399_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na873_1), .IN8(na3421_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a872_2 ( .OUT(na872_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na872_1_i) );
// C_MX2b/D///      x42y51     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a873_1 ( .OUT(na873_1_i), .IN1(na399_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na874_1), .IN8(na3420_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a873_2 ( .OUT(na873_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na873_1_i) );
// C_MX2a/D///      x40y53     80'h00_FE00_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a874_1 ( .OUT(na874_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na3417_1), .IN4(na875_1), .IN5(~na399_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a874_2 ( .OUT(na874_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na874_1_i) );
// C_MX2b/D///      x42y54     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a875_1 ( .OUT(na875_1_i), .IN1(~na399_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3416_2), .IN8(na876_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a875_2 ( .OUT(na875_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na875_1_i) );
// C_MX2a/D///      x38y54     80'h00_FE00_00_0040_0C0C_FA00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a876_1 ( .OUT(na876_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na397_1), .IN4(na3414_1), .IN5(na399_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a876_2 ( .OUT(na876_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na876_1_i) );
// C_MX4b////D      x23y63     80'h00_FA18_00_0040_0AF4_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a877_1 ( .OUT(na877_1), .IN1(1'b1), .IN2(na878_1), .IN3(1'b1), .IN4(~na864_1), .IN5(na1488_1), .IN6(na4301_2), .IN7(~na880_2),
                     .IN8(na4443_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a877_5 ( .OUT(na877_2), .CLK(na1739_1), .EN(na1487_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na877_1) );
// C_MX2b////      x21y52     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a878_1 ( .OUT(na878_1), .IN1(~na2479_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4300_2), .IN8(na3256_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y40     80'h00_0018_00_0040_0A55_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a879_1 ( .OUT(na879_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na203_2), .IN5(~na698_1), .IN6(1'b0), .IN7(~na3532_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x26y59     80'h00_0060_00_0000_0C08_FFCB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a880_4 ( .OUT(na880_2), .IN1(na3585_1), .IN2(~na2474_1), .IN3(1'b0), .IN4(na214_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////D      x35y52     80'h00_FA18_00_0000_0666_F3B5
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a881_1 ( .OUT(na881_1), .IN1(na882_2), .IN2(1'b1), .IN3(~na3588_1), .IN4(na864_1), .IN5(1'b1), .IN6(na1482_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a881_5 ( .OUT(na881_2), .CLK(na1739_1), .EN(na1481_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na881_1) );
// C_///AND/      x19y59     80'h00_0060_00_0000_0C08_FF31
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a882_4 ( .OUT(na882_2), .IN1(~na883_1), .IN2(~na2478_1), .IN3(1'b1), .IN4(~na3256_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x19y57     80'h00_0018_00_0000_0888_F9AC
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a883_1 ( .OUT(na883_1), .IN1(1'b0), .IN2(~na4303_2), .IN3(~na2481_2), .IN4(1'b0), .IN5(na4524_2), .IN6(na2478_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x16y64     80'h00_0060_00_0000_0C08_FF2C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a884_4 ( .OUT(na884_2), .IN1(1'b1), .IN2(na4119_2), .IN3(na1369_1), .IN4(~na214_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x20y52     80'h00_0018_00_0000_0C88_DCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a885_1 ( .OUT(na885_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na4297_2), .IN7(~na2481_2), .IN8(na3589_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x25y59     80'h00_F600_00_0040_0C0A_2F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a886_1 ( .OUT(na886_1_i), .IN1(1'b0), .IN2(na881_1), .IN3(1'b0), .IN4(na2499_1), .IN5(1'b1), .IN6(1'b1), .IN7(na304_1), .IN8(~na4164_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a886_2 ( .OUT(na886_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na886_1_i) );
// C_///AND/D      x24y51     80'h00_FE00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a887_4 ( .OUT(na887_2_i), .IN1(na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(na3426_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a887_5 ( .OUT(na887_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na887_2_i) );
// C_AND////D      x23y57     80'h00_FE18_00_0000_0888_33FC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a888_1 ( .OUT(na888_1), .IN1(1'b1), .IN2(na927_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na927_1), .IN7(1'b1), .IN8(~na1303_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a888_5 ( .OUT(na888_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na888_1) );
// C_ANDXOR/D//AND/D      x16y49     80'h00_FA00_80_0000_0C68_CEAF
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a891_1 ( .OUT(na891_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na3590_1), .IN6(~na2474_2), .IN7(1'b1), .IN8(~na4299_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a891_2 ( .OUT(na891_1), .CLK(na1739_1), .EN(na1479_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na891_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a891_4 ( .OUT(na891_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na891_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a891_5 ( .OUT(na891_2), .CLK(na1739_1), .EN(na1479_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na891_2_i) );
// C_ORAND*/D//ORAND*/D      x46y49     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a892_1 ( .OUT(na892_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na4305_2), .IN7(~na2593_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a892_2 ( .OUT(na892_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na892_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a892_4 ( .OUT(na892_2_i), .IN1(~na301_1), .IN2(~na894_1), .IN3(~na2593_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a892_5 ( .OUT(na892_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na892_2_i) );
// C_ORAND*/D//ORAND*/D      x43y50     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a894_1 ( .OUT(na894_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na894_2), .IN7(~na2595_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a894_2 ( .OUT(na894_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na894_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a894_4 ( .OUT(na894_2_i), .IN1(~na301_1), .IN2(~na4308_2), .IN3(~na2595_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a894_5 ( .OUT(na894_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na894_2_i) );
// C_ORAND*/D//ORAND*/D      x46y50     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a896_1 ( .OUT(na896_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na4309_2), .IN7(~na2597_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a896_2 ( .OUT(na896_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na896_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a896_4 ( .OUT(na896_2_i), .IN1(~na301_1), .IN2(~na898_1), .IN3(~na2597_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a896_5 ( .OUT(na896_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na896_2_i) );
// C_ORAND*/D//ORAND*/D      x39y50     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a898_1 ( .OUT(na898_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na898_2), .IN7(~na2599_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a898_2 ( .OUT(na898_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na898_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a898_4 ( .OUT(na898_2_i), .IN1(~na301_1), .IN2(~na900_1), .IN3(~na2599_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a898_5 ( .OUT(na898_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na898_2_i) );
// C_ORAND*/D//ORAND*/D      x41y50     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a900_1 ( .OUT(na900_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na900_2), .IN7(~na1819_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a900_2 ( .OUT(na900_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na900_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a900_4 ( .OUT(na900_2_i), .IN1(~na301_1), .IN2(~na902_1), .IN3(~na1819_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a900_5 ( .OUT(na900_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na900_2_i) );
// C_ORAND*/D//ORAND*/D      x41y46     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a902_1 ( .OUT(na902_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na902_2), .IN7(~na1821_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a902_2 ( .OUT(na902_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na902_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a902_4 ( .OUT(na902_2_i), .IN1(~na301_1), .IN2(~na904_1), .IN3(~na1821_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a902_5 ( .OUT(na902_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na902_2_i) );
// C_ORAND*/D//ORAND*/D      x45y48     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a904_1 ( .OUT(na904_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na904_2), .IN7(~na1823_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a904_2 ( .OUT(na904_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na904_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a904_4 ( .OUT(na904_2_i), .IN1(~na301_1), .IN2(~na906_1), .IN3(~na1823_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a904_5 ( .OUT(na904_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na904_2_i) );
// C_ORAND*/D//ORAND*/D      x41y48     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a906_1 ( .OUT(na906_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na906_2), .IN7(~na1825_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a906_2 ( .OUT(na906_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na906_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a906_4 ( .OUT(na906_2_i), .IN1(~na301_1), .IN2(~na4318_2), .IN3(~na1825_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a906_5 ( .OUT(na906_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na906_2_i) );
// C_ORAND*/D//ORAND*/D      x45y47     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a908_1 ( .OUT(na908_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na4319_2), .IN7(~na1811_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a908_2 ( .OUT(na908_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na908_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a908_4 ( .OUT(na908_2_i), .IN1(~na301_1), .IN2(~na910_1), .IN3(~na1811_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a908_5 ( .OUT(na908_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na908_2_i) );
// C_ORAND*/D//ORAND*/D      x47y46     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a910_1 ( .OUT(na910_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na910_2), .IN7(~na1813_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a910_2 ( .OUT(na910_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na910_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a910_4 ( .OUT(na910_2_i), .IN1(~na301_1), .IN2(~na912_1), .IN3(~na1813_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a910_5 ( .OUT(na910_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na910_2_i) );
// C_ORAND*/D//ORAND*/D      x43y46     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a912_1 ( .OUT(na912_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na912_2), .IN7(~na1815_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a912_2 ( .OUT(na912_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na912_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a912_4 ( .OUT(na912_2_i), .IN1(~na301_1), .IN2(~na914_1), .IN3(~na1815_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a912_5 ( .OUT(na912_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na912_2_i) );
// C_ORAND*/D//ORAND*/D      x45y46     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a914_1 ( .OUT(na914_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na914_2), .IN7(~na1817_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a914_2 ( .OUT(na914_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na914_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a914_4 ( .OUT(na914_2_i), .IN1(~na301_1), .IN2(~na916_1), .IN3(~na1817_1), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a914_5 ( .OUT(na914_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na914_2_i) );
// C_ORAND*/D//ORAND*/D      x45y42     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a916_1 ( .OUT(na916_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na916_2), .IN7(~na3532_1),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a916_2 ( .OUT(na916_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na916_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a916_4 ( .OUT(na916_2_i), .IN1(~na301_1), .IN2(~na4324_2), .IN3(~na3531_2), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a916_5 ( .OUT(na916_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na916_2_i) );
// C_ORAND*/D//ORAND*/D      x46y41     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a918_1 ( .OUT(na918_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na4325_2), .IN7(~na4608_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a918_2 ( .OUT(na918_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na918_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a918_4 ( .OUT(na918_2_i), .IN1(~na301_1), .IN2(~na920_1), .IN3(~na4607_2), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a918_5 ( .OUT(na918_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na918_2_i) );
// C_ORAND*/D//ORAND*/D      x43y42     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a920_1 ( .OUT(na920_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na920_2), .IN7(~na3528_1),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a920_2 ( .OUT(na920_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na920_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a920_4 ( .OUT(na920_2_i), .IN1(~na301_1), .IN2(~na4328_2), .IN3(~na3527_2), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a920_5 ( .OUT(na920_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na920_2_i) );
// C_ORAND*/D//ORAND*/D      x40y41     80'h00_F600_80_0000_0387_777D
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a922_1 ( .OUT(na922_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na301_1), .IN6(~na4329_2), .IN7(~na4606_2),
                     .IN8(~na302_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a922_2 ( .OUT(na922_1), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na922_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a922_4 ( .OUT(na922_2_i), .IN1(~na301_1), .IN2(na879_1), .IN3(~na4605_2), .IN4(~na302_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a922_5 ( .OUT(na922_2), .CLK(na1739_1), .EN(~na1404_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                     .D_IN(na922_2_i) );
// C_ORAND////      x33y53     80'h00_0018_00_0000_0C88_E3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a924_1 ( .OUT(na924_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na2474_1), .IN7(na4133_2), .IN8(na3657_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x26y70     80'h00_FE00_00_0040_0AC8_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a926_1 ( .OUT(na926_1_i), .IN1(1'b1), .IN2(na978_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4330_2),
                     .IN8(~na926_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a926_2 ( .OUT(na926_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na926_1_i) );
// C_AND/D//AND/D      x17y62     80'h00_FE00_80_0000_0C88_A5F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a927_1 ( .OUT(na927_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na436_1), .IN6(1'b1), .IN7(na1653_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a927_2 ( .OUT(na927_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na927_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a927_4 ( .OUT(na927_2_i), .IN1(~na436_1), .IN2(~na927_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a927_5 ( .OUT(na927_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na927_2_i) );
// C_MX4b/D///      x26y71     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a928_1 ( .OUT(na928_1_i), .IN1(1'b1), .IN2(~na978_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1658_1), .IN6(na4332_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a928_2 ( .OUT(na928_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na928_1_i) );
// C_MX4b/D///      x27y72     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a929_1 ( .OUT(na929_1_i), .IN1(1'b1), .IN2(~na978_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1658_2), .IN6(na929_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a929_2 ( .OUT(na929_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na929_1_i) );
// C_///OR/D      x13y47     80'h00_FE00_80_0000_0C0E_FFA5
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a930_4 ( .OUT(na930_2_i), .IN1(~na3259_1), .IN2(1'b0), .IN3(na931_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a930_5 ( .OUT(na930_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na930_2_i) );
// C_AND////      x22y53     80'h00_0018_00_0000_0888_32F2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a931_1 ( .OUT(na931_1), .IN1(na2479_2), .IN2(~na122_2), .IN3(1'b1), .IN4(1'b1), .IN5(na3218_1), .IN6(~na122_1), .IN7(1'b1),
                     .IN8(~na1495_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x21y44     80'h00_FE00_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a932_1 ( .OUT(na932_1_i), .IN1(1'b1), .IN2(na194_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na211_1), .IN8(na1545_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a932_2 ( .OUT(na932_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na932_1_i) );
// C_MX2b/D///      x23y42     80'h00_FE00_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a933_1 ( .OUT(na933_1_i), .IN1(1'b1), .IN2(na194_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4414_2), .IN8(na1545_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a933_2 ( .OUT(na933_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na933_1_i) );
// C_ORAND/D///      x20y37     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a934_1 ( .OUT(na934_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3661_1), .IN6(~na194_1), .IN7(~na3660_2),
                     .IN8(~na4536_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a934_2 ( .OUT(na934_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na934_1_i) );
// C_///ORAND/D      x20y35     80'h00_FE00_80_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a936_4 ( .OUT(na936_2_i), .IN1(~na3664_1), .IN2(~na194_1), .IN3(~na3660_2), .IN4(~na4537_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a936_5 ( .OUT(na936_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na936_2_i) );
// C_ORAND/D///      x19y36     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a938_1 ( .OUT(na938_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3667_1), .IN6(~na194_1), .IN7(~na3660_2),
                     .IN8(~na2489_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a938_2 ( .OUT(na938_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na938_1_i) );
// C_///ORAND/D      x19y36     80'h00_FE00_80_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a940_4 ( .OUT(na940_2_i), .IN1(~na3670_1), .IN2(~na194_1), .IN3(~na3660_2), .IN4(~na4538_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a940_5 ( .OUT(na940_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na940_2_i) );
// C_ORAND/D///      x20y35     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a942_1 ( .OUT(na942_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3673_1), .IN6(~na194_1), .IN7(~na3660_2),
                     .IN8(~na2489_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a942_2 ( .OUT(na942_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na942_1_i) );
// C_MX2b/D///      x42y41     80'h00_FE00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a944_1 ( .OUT(na944_1_i), .IN1(1'b1), .IN2(~na194_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3187_1), .IN6(na3674_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a944_2 ( .OUT(na944_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na944_1_i) );
// C_MX2b/D///      x39y37     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a945_1 ( .OUT(na945_1_i), .IN1(1'b1), .IN2(na194_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3675_1), .IN6(na3188_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a945_2 ( .OUT(na945_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na945_1_i) );
// C_MX2b/D///      x38y37     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a946_1 ( .OUT(na946_1_i), .IN1(1'b1), .IN2(na194_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3676_1), .IN6(na3189_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a946_2 ( .OUT(na946_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na946_1_i) );
// C_MX2b/D///      x40y37     80'h00_FE00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a947_1 ( .OUT(na947_1_i), .IN1(1'b1), .IN2(na194_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3677_1), .IN8(na3190_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a947_2 ( .OUT(na947_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na947_1_i) );
// C_MX2b/D///      x38y42     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a948_1 ( .OUT(na948_1_i), .IN1(1'b1), .IN2(na194_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3678_2), .IN6(na3191_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a948_2 ( .OUT(na948_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na948_1_i) );
// C_MX2b/D///      x39y41     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a949_1 ( .OUT(na949_1_i), .IN1(1'b1), .IN2(na194_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3679_1), .IN6(na3192_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a949_2 ( .OUT(na949_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na949_1_i) );
// C_MX2b/D///      x33y42     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a950_1 ( .OUT(na950_1_i), .IN1(1'b1), .IN2(na194_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3680_1), .IN6(na3193_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a950_2 ( .OUT(na950_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na950_1_i) );
// C_ORAND*////D      x22y59     80'h00_FE18_00_0000_0788_5BD3
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a951_1 ( .OUT(na951_1), .IN1(1'b0), .IN2(~na957_1), .IN3(~na304_1), .IN4(na3682_1), .IN5(na959_1), .IN6(~na957_2), .IN7(~na304_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a951_5 ( .OUT(na951_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na951_1) );
// C_AND///AND/      x26y61     80'h00_0078_00_0000_0C88_12C3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a952_1 ( .OUT(na952_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3683_1), .IN6(~na2474_1), .IN7(~na4523_2),
                     .IN8(~na2473_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a952_4 ( .OUT(na952_2), .IN1(1'b1), .IN2(~na2474_1), .IN3(1'b1), .IN4(na2473_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x17y54     80'h00_0060_00_0000_0C06_FFB3
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a953_4 ( .OUT(na953_2), .IN1(1'b1), .IN2(na878_1), .IN3(~na4611_2), .IN4(na954_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x22y50     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a954_1 ( .OUT(na954_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2472_1), .IN6(na4531_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x19y58     80'h00_0078_00_0000_0C88_8C51
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a957_1 ( .OUT(na957_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3258_2), .IN7(na123_1), .IN8(na3252_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a957_4 ( .OUT(na957_2), .IN1(~na4528_2), .IN2(~na2478_1), .IN3(~na2481_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y51     80'h00_0018_00_0040_0A33_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a959_1 ( .OUT(na959_1), .IN1(~na924_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(~na3688_2), .IN6(~na1593_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x21y54     80'h00_0060_00_0000_0C06_FFAC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a963_4 ( .OUT(na963_2), .IN1(1'b0), .IN2(na193_2), .IN3(na4523_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x27y59     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a964_1 ( .OUT(na964_1), .IN1(1'b1), .IN2(na2474_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3185_1), .IN8(na3186_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x33y43     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a965_1 ( .OUT(na965_1_i), .IN1(1'b1), .IN2(na194_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3694_2), .IN6(na3194_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a965_2 ( .OUT(na965_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na965_1_i) );
// C_MX2b////      x40y40     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a966_1 ( .OUT(na966_1), .IN1(1'b1), .IN2(na194_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4127_2), .IN8(na1545_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x39y40     80'h00_0018_00_0040_0AC4_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a967_1 ( .OUT(na967_1), .IN1(1'b1), .IN2(na194_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na4126_2), .IN8(na1545_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x25y42     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a968_4 ( .OUT(na968_2), .IN1(~na3661_1), .IN2(~na194_1), .IN3(~na969_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x26y45     80'h00_0018_00_0040_0AA0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a969_1 ( .OUT(na969_1), .IN1(1'b1), .IN2(~na194_1), .IN3(1'b1), .IN4(~na203_1), .IN5(1'b0), .IN6(na2482_1), .IN7(1'b0), .IN8(na853_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x22y46     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a970_4 ( .OUT(na970_2), .IN1(~na3664_1), .IN2(~na194_1), .IN3(~na971_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x26y43     80'h00_0018_00_0040_0AC0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a971_1 ( .OUT(na971_1), .IN1(1'b1), .IN2(na4124_2), .IN3(1'b1), .IN4(~na4122_2), .IN5(1'b0), .IN6(1'b0), .IN7(na856_1), .IN8(na2483_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x24y43     80'h00_0060_00_0000_0C08_FF37
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a972_4 ( .OUT(na972_2), .IN1(~na3667_1), .IN2(~na194_1), .IN3(1'b0), .IN4(~na973_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x26y44     80'h00_0018_00_0040_0A50_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a973_1 ( .OUT(na973_1), .IN1(1'b1), .IN2(na194_1), .IN3(1'b1), .IN4(na203_1), .IN5(na858_1), .IN6(1'b0), .IN7(na2484_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x25y42     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a974_1 ( .OUT(na974_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3670_1), .IN6(~na194_1), .IN7(~na975_1),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x30y45     80'h00_0018_00_0040_0AA0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a975_1 ( .OUT(na975_1), .IN1(1'b1), .IN2(~na194_1), .IN3(1'b1), .IN4(~na203_1), .IN5(1'b0), .IN6(na2485_2), .IN7(1'b0), .IN8(na860_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x25y41     80'h00_0060_00_0000_0C08_FF37
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a976_4 ( .OUT(na976_2), .IN1(~na3673_1), .IN2(~na194_1), .IN3(1'b0), .IN4(~na977_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x26y42     80'h00_0018_00_0040_0AA0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a977_1 ( .OUT(na977_1), .IN1(1'b1), .IN2(~na194_1), .IN3(1'b1), .IN4(~na203_1), .IN5(1'b0), .IN6(na2486_1), .IN7(1'b0), .IN8(na862_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x27y70     80'h00_FE00_00_0000_0C88_CEFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a978_1 ( .OUT(na978_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na445_2), .IN6(na978_1), .IN7(1'b0), .IN8(na3695_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a978_2 ( .OUT(na978_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na978_1_i) );
// C_///AND/D      x62y87     80'h00_FE00_80_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a980_4 ( .OUT(na980_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1149_2), .IN4(na1649_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a980_5 ( .OUT(na980_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na980_2_i) );
// C_///AND/      x36y69     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a982_4 ( .OUT(na982_2), .IN1(na408_1), .IN2(1'b1), .IN3(~na407_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y71     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a983_4 ( .OUT(na983_2), .IN1(~na7_2), .IN2(1'b1), .IN3(na11_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x31y73     80'h00_FE00_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a984_1 ( .OUT(na984_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3698_1), .IN6(~na3697_2), .IN7(~na1149_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a984_2 ( .OUT(na984_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na984_1_i) );
// C_AND/D//AND/D      x56y92     80'h00_FE00_80_0000_0C88_2F4F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a986_1 ( .OUT(na986_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1651_1), .IN8(~na4366_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a986_2 ( .OUT(na986_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na986_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a986_4 ( .OUT(na986_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na1149_2), .IN4(na1649_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a986_5 ( .OUT(na986_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na986_2_i) );
// C_AND/D///      x59y69     80'h00_FE00_00_0000_0888_8141
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a987_1 ( .OUT(na987_1_i), .IN1(~na4423_2), .IN2(~na285_2), .IN3(~na1149_2), .IN4(na4153_2), .IN5(~na987_1), .IN6(~na22_2),
                     .IN7(na4070_2), .IN8(na4111_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a987_2 ( .OUT(na987_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na987_1_i) );
// C_AND////      x20y89     80'h00_0018_00_0000_0888_1125
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a990_1 ( .OUT(na990_1), .IN1(~na411_1), .IN2(1'b1), .IN3(na992_1), .IN4(~na413_1), .IN5(~na418_1), .IN6(~na412_1), .IN7(~na1351_2),
                     .IN8(~na1350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x22y81     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a992_1 ( .OUT(na992_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na414_1), .IN6(~na415_1), .IN7(~na416_1), .IN8(~na417_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x40y78     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a993_1 ( .OUT(na993_1_i), .IN1(~na399_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3424_1), .IN8(na994_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a993_2 ( .OUT(na993_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na993_1_i) );
// C_MX2b/D///      x38y60     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a994_1 ( .OUT(na994_1_i), .IN1(~na399_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3423_2), .IN8(na995_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a994_2 ( .OUT(na994_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na994_1_i) );
// C_MX2b/D///      x38y56     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a995_1 ( .OUT(na995_1_i), .IN1(na399_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na996_1), .IN8(na3421_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a995_2 ( .OUT(na995_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na995_1_i) );
// C_MX2b/D///      x40y51     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a996_1 ( .OUT(na996_1_i), .IN1(na399_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na997_1), .IN8(na3420_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a996_2 ( .OUT(na996_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na996_1_i) );
// C_MX2b/D///      x36y53     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a997_1 ( .OUT(na997_1_i), .IN1(~na399_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3417_1), .IN8(na998_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a997_2 ( .OUT(na997_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na997_1_i) );
// C_MX2b/D///      x34y54     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a998_1 ( .OUT(na998_1_i), .IN1(~na399_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3416_2), .IN8(na999_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a998_2 ( .OUT(na998_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na998_1_i) );
// C_MX2b/D///      x40y54     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a999_1 ( .OUT(na999_1_i), .IN1(na399_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na398_1), .IN8(na3414_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a999_2 ( .OUT(na999_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na999_1_i) );
// C_MX2b/D///      x39y75     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1000_1 ( .OUT(na1000_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1001_1), .IN8(na2846_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1000_2 ( .OUT(na1000_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1000_1_i) );
// C_MX2b/D///      x42y79     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1001_1 ( .OUT(na1001_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1002_1), .IN8(na1780_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1001_2 ( .OUT(na1001_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1001_1_i) );
// C_MX2b/D///      x44y79     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1002_1 ( .OUT(na1002_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1003_1), .IN8(na1780_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1002_2 ( .OUT(na1002_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1002_1_i) );
// C_MX2b/D///      x42y77     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1003_1 ( .OUT(na1003_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1004_1), .IN8(na1782_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1003_2 ( .OUT(na1003_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1003_1_i) );
// C_MX2b/D///      x40y71     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1004_1 ( .OUT(na1004_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4335_2), .IN8(na1782_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1004_2 ( .OUT(na1004_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1004_1_i) );
// C_MX2b/D///      x43y82     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1005_1 ( .OUT(na1005_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1006_1), .IN8(na1792_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1005_2 ( .OUT(na1005_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1005_1_i) );
// C_MX2b/D///      x44y81     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1006_1 ( .OUT(na1006_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1007_1), .IN8(na1792_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1006_2 ( .OUT(na1006_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1006_1_i) );
// C_MX2b/D///      x46y77     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1007_1 ( .OUT(na1007_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1008_1), .IN8(na1794_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1007_2 ( .OUT(na1007_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1007_1_i) );
// C_MX2b/D///      x44y73     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1008_1 ( .OUT(na1008_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1009_1), .IN8(na1794_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1008_2 ( .OUT(na1008_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1008_1_i) );
// C_MX2b/D///      x40y65     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1009_1 ( .OUT(na1009_1_i), .IN1(1'b1), .IN2(na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3424_1), .IN8(na1010_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1009_2 ( .OUT(na1009_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1009_1_i) );
// C_MX2b/D///      x40y66     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1010_1 ( .OUT(na1010_1_i), .IN1(1'b1), .IN2(na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3423_2), .IN8(na1011_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1010_2 ( .OUT(na1010_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1010_1_i) );
// C_MX2b/D///      x40y60     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1011_1 ( .OUT(na1011_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1012_1), .IN8(na3421_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1011_2 ( .OUT(na1011_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1011_1_i) );
// C_MX2b/D///      x38y59     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1012_1 ( .OUT(na1012_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1013_1), .IN8(na3420_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1012_2 ( .OUT(na1012_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1012_1_i) );
// C_MX2b/D///      x36y61     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1013_1 ( .OUT(na1013_1_i), .IN1(1'b1), .IN2(na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3417_1), .IN8(na1014_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1013_2 ( .OUT(na1013_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1013_1_i) );
// C_MX2b/D///      x36y66     80'h00_F600_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1014_1 ( .OUT(na1014_1_i), .IN1(1'b1), .IN2(na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3416_2), .IN8(na1597_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1014_2 ( .OUT(na1014_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1014_1_i) );
// C_MX2b/D///      x40y75     80'h00_F600_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1015_1 ( .OUT(na1015_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2714_1), .IN6(na4562_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1015_2 ( .OUT(na1015_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1015_1_i) );
// C_MX2b/D///      x41y82     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1016_1 ( .OUT(na1016_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1017_1), .IN8(na1792_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1016_2 ( .OUT(na1016_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1016_1_i) );
// C_MX2b/D///      x42y81     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1017_1 ( .OUT(na1017_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1018_1), .IN8(na1784_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1017_2 ( .OUT(na1017_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1017_1_i) );
// C_MX2b/D///      x40y79     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1018_1 ( .OUT(na1018_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1019_1), .IN8(na1784_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1018_2 ( .OUT(na1018_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1018_1_i) );
// C_MX2b/D///      x50y87     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1019_1 ( .OUT(na1019_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1020_1), .IN8(na1786_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1019_2 ( .OUT(na1019_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1019_1_i) );
// C_MX2b/D///      x46y81     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1020_1 ( .OUT(na1020_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1021_1), .IN8(na1786_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1020_2 ( .OUT(na1020_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1020_1_i) );
// C_MX2b/D///      x48y81     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1021_1 ( .OUT(na1021_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1022_1), .IN8(na1788_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1021_2 ( .OUT(na1021_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1021_1_i) );
// C_MX2b/D///      x44y77     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1022_1 ( .OUT(na1022_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1023_1), .IN8(na1788_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1022_2 ( .OUT(na1022_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1022_1_i) );
// C_MX2b/D///      x48y77     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1023_1 ( .OUT(na1023_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1024_1), .IN8(na1790_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1023_2 ( .OUT(na1023_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1023_1_i) );
// C_MX2b/D///      x40y77     80'h00_F600_00_0040_0AC4_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1024_1 ( .OUT(na1024_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1025_1), .IN8(na1790_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1024_2 ( .OUT(na1024_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1024_1_i) );
// C_MX2b////      x38y75     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1025_1 ( .OUT(na1025_1), .IN1(1'b1), .IN2(~na4551_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2714_1), .IN6(~na1005_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x50y85     80'h00_FE00_00_0040_0C0A_3F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1026_1 ( .OUT(na1026_1_i), .IN1(1'b0), .IN2(na1029_1), .IN3(1'b0), .IN4(na1027_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1028_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1026_2 ( .OUT(na1026_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1026_1_i) );
// C_MX2b////      x48y82     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1027_1 ( .OUT(na1027_1), .IN1(na218_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1026_1), .IN8(na1786_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y86     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1028_1 ( .OUT(na1028_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2712_2), .IN6(na232_1), .IN7(na2713_1), .IN8(na2707_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x47y82     80'h00_FE00_00_0040_0C05_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1029_1 ( .OUT(na1029_1_i), .IN1(na1030_1), .IN2(1'b0), .IN3(na1031_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1028_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1029_2 ( .OUT(na1029_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1029_1_i) );
// C_MX2b////      x49y79     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1030_1 ( .OUT(na1030_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4135_2), .IN5(1'b0), .IN6(na1029_1), .IN7(1'b0), .IN8(na1788_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x50y81     80'h00_FE00_00_0040_0C05_C000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1031_1 ( .OUT(na1031_1_i), .IN1(na1032_1), .IN2(1'b0), .IN3(na1033_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1028_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1031_2 ( .OUT(na1031_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1031_1_i) );
// C_MX2b////      x49y81     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1032_1 ( .OUT(na1032_1), .IN1(na218_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1031_1), .IN8(na1788_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x48y83     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1033_1 ( .OUT(na1033_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1028_1), .IN5(na1034_1), .IN6(1'b0), .IN7(na1035_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1033_2 ( .OUT(na1033_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1033_1_i) );
// C_MX2b////      x47y77     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1034_1 ( .OUT(na1034_1), .IN1(na218_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1033_1), .IN8(na1790_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x48y79     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1035_1 ( .OUT(na1035_1_i), .IN1(na218_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1028_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1035_1),
                      .IN8(na1790_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1035_2 ( .OUT(na1035_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1035_1_i) );
// C_MX4b/D///      x35y75     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1036_1 ( .OUT(na1036_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1036_1), .IN6(na66_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1036_2 ( .OUT(na1036_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1036_1_i) );
// C_MX4b////D      x39y89     80'h00_FA18_00_0040_0AF4_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1037_1 ( .OUT(na1037_1), .IN1(1'b1), .IN2(na4338_2), .IN3(1'b1), .IN4(~na993_1), .IN5(na1510_1), .IN6(na4339_2), .IN7(~na1043_1),
                      .IN8(na4450_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1037_5 ( .OUT(na1037_2), .CLK(na1739_1), .EN(na232_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1037_1) );
// C_MX2a////      x36y85     80'h00_0018_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1038_1 ( .OUT(na1038_1), .IN1(na1042_1), .IN2(na3701_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na2712_1), .IN6(1'b1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x40y80     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1039_1 ( .OUT(na1039_1), .IN1(~na1040_2), .IN2(1'b1), .IN3(na4141_2), .IN4(1'b1), .IN5(na1000_1), .IN6(na1005_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x45y83     80'h00_0060_00_0000_0C08_FF12
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1040_4 ( .OUT(na1040_2), .IN1(na2712_1), .IN2(~na4550_2), .IN3(~na2713_2), .IN4(~na2710_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x41y63     80'h00_0018_00_0040_0ACC_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1042_1 ( .OUT(na1042_1), .IN1(~na399_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na3424_1), .IN8(~na871_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x42y89     80'h00_0018_00_0000_0C88_BCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1043_1 ( .OUT(na1043_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na232_2), .IN7(na3703_1), .IN8(~na2707_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////D      x49y92     80'h00_FA18_00_0000_0666_F3B5
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1044_1 ( .OUT(na1044_1), .IN1(na1045_2), .IN2(1'b1), .IN3(~na3706_1), .IN4(na993_1), .IN5(1'b1), .IN6(na1504_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1044_5 ( .OUT(na1044_2), .CLK(na1739_1), .EN(na1503_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1044_1) );
// C_///AND/      x49y87     80'h00_0060_00_0000_0C08_FF31
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1045_4 ( .OUT(na1045_2), .IN1(~na2712_2), .IN2(~na3701_2), .IN3(1'b1), .IN4(~na1046_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x38y88     80'h00_0018_00_0000_0888_9FAC
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1046_1 ( .OUT(na1046_1), .IN1(1'b0), .IN2(~na1047_1), .IN3(~na2713_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2713_2),
                      .IN8(na2710_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y92     80'h00_0018_00_0000_0C88_4CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1047_1 ( .OUT(na1047_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1048_1), .IN7(~na432_2), .IN8(na239_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x33y92     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1048_1 ( .OUT(na1048_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na434_2), .IN6(1'b1), .IN7(~na4199_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x40y84     80'h00_0018_00_0000_0C88_DCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1049_1 ( .OUT(na1049_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na4334_2), .IN7(~na2713_1), .IN8(na3707_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x48y92     80'h00_F600_00_0040_0C0A_2F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1050_1 ( .OUT(na1050_1_i), .IN1(1'b0), .IN2(na1044_1), .IN3(1'b0), .IN4(na2739_1), .IN5(1'b1), .IN6(1'b1), .IN7(na226_1),
                      .IN8(~na1347_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1050_2 ( .OUT(na1050_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1050_1_i) );
// C_ANDXOR/D//AND/D      x29y92     80'h00_FA00_80_0000_0C68_EAFC
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1051_1 ( .OUT(na1051_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na4337_2), .IN6(1'b1), .IN7(~na3708_2),
                      .IN8(~na2707_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1051_2 ( .OUT(na1051_1), .CLK(na1739_1), .EN(na1501_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1051_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1051_4 ( .OUT(na1051_2_i), .IN1(1'b1), .IN2(na1051_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1051_5 ( .OUT(na1051_2), .CLK(na1739_1), .EN(na1501_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1051_2_i) );
// C_ORAND*/D//ORAND*/D      x59y72     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1052_1 ( .OUT(na1052_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4341_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na2840_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1052_2 ( .OUT(na1052_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1052_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1052_4 ( .OUT(na1052_2_i), .IN1(~na1054_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na2840_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1052_5 ( .OUT(na1052_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1052_2_i) );
// C_ORAND*/D//ORAND*/D      x57y71     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1054_1 ( .OUT(na1054_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1054_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na2842_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1054_2 ( .OUT(na1054_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1054_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1054_4 ( .OUT(na1054_2_i), .IN1(~na1056_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na2842_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1054_5 ( .OUT(na1054_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1054_2_i) );
// C_ORAND*/D//ORAND*/D      x57y75     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1056_1 ( .OUT(na1056_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1056_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na2844_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1056_2 ( .OUT(na1056_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1056_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1056_4 ( .OUT(na1056_2_i), .IN1(~na4342_2), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na2844_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1056_5 ( .OUT(na1056_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1056_2_i) );
// C_ORAND*/D//ORAND*/D      x56y75     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1058_1 ( .OUT(na1058_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4343_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na2846_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1058_2 ( .OUT(na1058_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1058_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1058_4 ( .OUT(na1058_2_i), .IN1(~na1060_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na2846_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1058_5 ( .OUT(na1058_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1058_2_i) );
// C_ORAND*/D//ORAND*/D      x57y79     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1060_1 ( .OUT(na1060_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1060_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na1780_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1060_2 ( .OUT(na1060_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1060_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1060_4 ( .OUT(na1060_2_i), .IN1(~na1062_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na1780_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1060_5 ( .OUT(na1060_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1060_2_i) );
// C_ORAND*/D//ORAND*/D      x55y79     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1062_1 ( .OUT(na1062_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1062_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na1782_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1062_2 ( .OUT(na1062_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1062_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1062_4 ( .OUT(na1062_2_i), .IN1(~na1064_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na1782_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1062_5 ( .OUT(na1062_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1062_2_i) );
// C_ORAND*/D//ORAND*/D      x55y81     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1064_1 ( .OUT(na1064_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1064_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na1784_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1064_2 ( .OUT(na1064_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1064_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1064_4 ( .OUT(na1064_2_i), .IN1(~na1066_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na1784_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1064_5 ( .OUT(na1064_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1064_2_i) );
// C_ORAND*/D//ORAND*/D      x53y81     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1066_1 ( .OUT(na1066_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1066_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na1786_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1066_2 ( .OUT(na1066_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1066_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1066_4 ( .OUT(na1066_2_i), .IN1(~na1068_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na1786_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1066_5 ( .OUT(na1066_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1066_2_i) );
// C_ORAND*/D//ORAND*/D      x61y79     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1068_1 ( .OUT(na1068_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1068_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na1788_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1068_2 ( .OUT(na1068_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1068_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1068_4 ( .OUT(na1068_2_i), .IN1(~na1070_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na1788_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1068_5 ( .OUT(na1068_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1068_2_i) );
// C_ORAND*/D//ORAND*/D      x59y79     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1070_1 ( .OUT(na1070_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1070_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na1790_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1070_2 ( .OUT(na1070_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1070_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1070_4 ( .OUT(na1070_2_i), .IN1(~na1072_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na1790_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1070_5 ( .OUT(na1070_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1070_2_i) );
// C_ORAND*/D//ORAND*/D      x57y81     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1072_1 ( .OUT(na1072_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1072_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na1792_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1072_2 ( .OUT(na1072_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1072_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1072_4 ( .OUT(na1072_2_i), .IN1(~na1074_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na1792_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1072_5 ( .OUT(na1072_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1072_2_i) );
// C_ORAND*/D//ORAND*/D      x57y77     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1074_1 ( .OUT(na1074_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1074_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na1794_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1074_2 ( .OUT(na1074_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1074_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1074_4 ( .OUT(na1074_2_i), .IN1(~na1076_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na1794_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1074_5 ( .OUT(na1074_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1074_2_i) );
// C_ORAND*/D//ORAND*/D      x55y71     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1076_1 ( .OUT(na1076_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1076_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na4594_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1076_2 ( .OUT(na1076_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1076_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1076_4 ( .OUT(na1076_2_i), .IN1(~na1078_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na4593_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1076_5 ( .OUT(na1076_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1076_2_i) );
// C_ORAND*/D//ORAND*/D      x55y69     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1078_1 ( .OUT(na1078_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1078_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na3421_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1078_2 ( .OUT(na1078_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1078_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1078_4 ( .OUT(na1078_2_i), .IN1(~na4361_2), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na3420_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1078_5 ( .OUT(na1078_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1078_2_i) );
// C_ORAND*/D//ORAND*/D      x56y72     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1080_1 ( .OUT(na1080_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4362_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na4592_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1080_2 ( .OUT(na1080_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1080_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1080_4 ( .OUT(na1080_2_i), .IN1(~na1082_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na4591_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1080_5 ( .OUT(na1080_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1080_2_i) );
// C_ORAND*/D//ORAND*/D      x51y71     80'h00_F600_80_0000_0387_777B
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1082_1 ( .OUT(na1082_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1082_2), .IN6(~na223_2), .IN7(~na224_1),
                      .IN8(~na3414_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1082_2 ( .OUT(na1082_1), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1082_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1082_4 ( .OUT(na1082_2_i), .IN1(na1042_1), .IN2(~na223_2), .IN3(~na224_1), .IN4(~na3413_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1082_5 ( .OUT(na1082_2), .CLK(na1739_1), .EN(~na1401_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1082_2_i) );
// C_///ORAND/      x60y87     80'h00_0060_00_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1084_4 ( .OUT(na1084_2), .IN1(na434_1), .IN2(na3775_2), .IN3(1'b0), .IN4(~na2707_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x58y82     80'h00_FE00_00_0000_0C88_5EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1085_1 ( .OUT(na1085_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1086_1), .IN6(na3777_2), .IN7(~na1149_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1085_2 ( .OUT(na1085_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1085_1_i) );
// C_MX4a////      x61y75     80'h00_0018_00_0040_0C82_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1086_1 ( .OUT(na1086_1), .IN1(1'b0), .IN2(na3778_1), .IN3(1'b0), .IN4(1'b1), .IN5(na1089_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1990_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x67y74     80'h00_0018_00_0040_0CCC_F100
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1087_1 ( .OUT(na1087_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na511_1), .IN4(~na1088_1), .IN5(~na4483_2), .IN6(~na1986_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x64y66     80'h00_0018_00_0000_0C88_C6FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1088_1 ( .OUT(na1088_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na535_1), .IN6(~na512_1), .IN7(1'b0), .IN8(~na1443_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x67y77     80'h00_0060_00_0000_0C08_FF28
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1089_4 ( .OUT(na1089_2), .IN1(na4101_2), .IN2(na1993_2), .IN3(na38_2), .IN4(~na1990_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x62y72     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1090_1 ( .OUT(na1090_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4101_2), .IN6(1'b1), .IN7(na38_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1090_2 ( .OUT(na1090_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1090_1_i) );
// C_///OR/D      x41y70     80'h00_FE00_80_0000_0C0E_FF0D
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1091_4 ( .OUT(na1091_2_i), .IN1(~na3578_1), .IN2(na1092_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1091_5 ( .OUT(na1091_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1091_2_i) );
// C_AND////      x43y86     80'h00_0018_00_0000_0888_53A2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1092_1 ( .OUT(na1092_1), .IN1(na2712_1), .IN2(~na819_2), .IN3(na3146_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na219_2), .IN7(~na1517_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x41y71     80'h00_FE00_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1093_1 ( .OUT(na1093_1_i), .IN1(1'b1), .IN2(na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na410_1), .IN6(na1543_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1093_2 ( .OUT(na1093_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1093_1_i) );
// C_MX2b/D///      x43y72     80'h00_FE00_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1094_1 ( .OUT(na1094_1_i), .IN1(1'b1), .IN2(na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na4197_2), .IN6(na1543_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1094_2 ( .OUT(na1094_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1094_1_i) );
// C_ORAND/D///      x37y68     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1095_1 ( .OUT(na1095_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3783_1), .IN6(~na817_1), .IN7(~na3782_1),
                      .IN8(~na2720_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1095_2 ( .OUT(na1095_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1095_1_i) );
// C_///ORAND/D      x39y68     80'h00_FE00_80_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1097_4 ( .OUT(na1097_2_i), .IN1(~na3786_1), .IN2(~na817_1), .IN3(~na3782_1), .IN4(~na2721_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1097_5 ( .OUT(na1097_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1097_2_i) );
// C_///ORAND/D      x39y65     80'h00_FE00_80_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1099_4 ( .OUT(na1099_2_i), .IN1(~na3789_1), .IN2(~na817_1), .IN3(~na3782_1), .IN4(~na2722_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1099_5 ( .OUT(na1099_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1099_2_i) );
// C_///ORAND/D      x37y68     80'h00_FE00_80_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1101_4 ( .OUT(na1101_2_i), .IN1(~na3792_1), .IN2(~na817_1), .IN3(~na3782_1), .IN4(~na2723_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1101_5 ( .OUT(na1101_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1101_2_i) );
// C_ORAND/D///      x35y59     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1103_1 ( .OUT(na1103_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3795_1), .IN6(~na817_1), .IN7(~na3782_1),
                      .IN8(~na2722_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1103_2 ( .OUT(na1103_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1103_1_i) );
// C_MX2b/D///      x49y68     80'h00_FE00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1105_1 ( .OUT(na1105_1_i), .IN1(1'b1), .IN2(~na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3199_1), .IN6(na3796_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1105_2 ( .OUT(na1105_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1105_1_i) );
// C_MX2b/D///      x49y65     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1106_1 ( .OUT(na1106_1_i), .IN1(1'b1), .IN2(~na817_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3200_1), .IN8(na3797_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1106_2 ( .OUT(na1106_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1106_1_i) );
// C_MX2b/D///      x50y67     80'h00_FE00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1107_1 ( .OUT(na1107_1_i), .IN1(1'b1), .IN2(na817_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3798_2), .IN8(na3201_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1107_2 ( .OUT(na1107_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1107_1_i) );
// C_MX2b/D///      x49y69     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1108_1 ( .OUT(na1108_1_i), .IN1(1'b1), .IN2(na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3799_2), .IN6(na3202_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1108_2 ( .OUT(na1108_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1108_1_i) );
// C_MX2b/D///      x45y68     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1109_1 ( .OUT(na1109_1_i), .IN1(1'b1), .IN2(na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3800_1), .IN6(na3203_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1109_2 ( .OUT(na1109_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1109_1_i) );
// C_MX2b/D///      x43y64     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1110_1 ( .OUT(na1110_1_i), .IN1(1'b1), .IN2(na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3801_1), .IN6(na3204_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1110_2 ( .OUT(na1110_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1110_1_i) );
// C_MX2b/D///      x46y69     80'h00_FE00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1111_1 ( .OUT(na1111_1_i), .IN1(1'b1), .IN2(na817_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3802_1), .IN8(na3205_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1111_2 ( .OUT(na1111_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1111_1_i) );
// C_ORAND*////D      x49y90     80'h00_FE18_00_0000_0788_5DD5
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1112_1 ( .OUT(na1112_1), .IN1(~na1118_1), .IN2(1'b0), .IN3(~na226_1), .IN4(na3804_1), .IN5(~na1118_2), .IN6(na1129_1), .IN7(~na226_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1112_5 ( .OUT(na1112_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1112_1) );
// C_AND///AND/      x44y92     80'h00_0078_00_0000_0C88_123C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1113_1 ( .OUT(na1113_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3805_2), .IN6(~na2706_1), .IN7(~na4548_2),
                      .IN8(~na2707_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1113_4 ( .OUT(na1113_2), .IN1(1'b1), .IN2(na2706_1), .IN3(1'b1), .IN4(~na2707_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x35y85     80'h00_0018_00_0000_0C66_5B00
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1114_1 ( .OUT(na1114_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na4613_2), .IN6(na1115_2), .IN7(na1038_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y76     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1115_4 ( .OUT(na1115_2), .IN1(na2712_1), .IN2(1'b1), .IN3(na2705_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x35y87     80'h00_0078_00_0000_0C88_8A51
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1118_1 ( .OUT(na1118_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3809_1), .IN6(1'b1), .IN7(na3815_2), .IN8(na1337_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1118_4 ( .OUT(na1118_2), .IN1(~na2712_2), .IN2(~na4553_2), .IN3(~na2713_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x33y89     80'h00_0060_00_0000_0C08_FFBA
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1120_4 ( .OUT(na1120_2), .IN1(na1292_1), .IN2(1'b0), .IN3(na3811_2), .IN4(~na1121_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x38y84     80'h00_0018_00_0040_0C61_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1121_1 ( .OUT(na1121_1), .IN1(na2712_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b0), .IN5(1'b1), .IN6(na4553_2), .IN7(1'b1), .IN8(na2710_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x38y91     80'h00_0060_00_0000_0C08_FFB5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1122_4 ( .OUT(na1122_2), .IN1(~na3812_1), .IN2(1'b0), .IN3(na3815_2), .IN4(~na2739_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x34y92     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1127_4 ( .OUT(na1127_2), .IN1(na1292_1), .IN2(na1506_1), .IN3(1'b0), .IN4(na1128_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x36y90     80'h00_0060_00_0000_0C08_FF4C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1128_4 ( .OUT(na1128_2), .IN1(1'b1), .IN2(na1048_1), .IN3(~na432_2), .IN4(na240_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x51y90     80'h00_0018_00_0040_0A55_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1129_1 ( .OUT(na1129_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na1084_2), .IN4(1'b1), .IN5(~na3816_2), .IN6(1'b0), .IN7(~na1599_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x37y91     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1133_1 ( .OUT(na1133_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na391_2), .IN7(1'b0), .IN8(na2707_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x41y89     80'h00_0018_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1134_1 ( .OUT(na1134_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2707_1), .IN5(1'b0), .IN6(na3197_1), .IN7(1'b0), .IN8(na3198_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x48y69     80'h00_FE00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1135_1 ( .OUT(na1135_1_i), .IN1(1'b1), .IN2(~na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3206_1), .IN6(na3822_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1135_2 ( .OUT(na1135_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1135_1_i) );
// C_MX2b////      x47y72     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1136_1 ( .OUT(na1136_1), .IN1(1'b1), .IN2(na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na4409_2), .IN6(na1543_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y71     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1137_1 ( .OUT(na1137_1), .IN1(1'b1), .IN2(na817_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na4408_2), .IN6(na1543_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x41y66     80'h00_0018_00_0000_0C88_37FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1138_1 ( .OUT(na1138_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3783_1), .IN6(~na817_1), .IN7(1'b0), .IN8(~na1139_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y74     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1139_1 ( .OUT(na1139_1), .IN1(na399_1), .IN2(1'b1), .IN3(~na4293_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1026_1),
                      .IN8(na2715_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x39y68     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1140_1 ( .OUT(na1140_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3786_1), .IN6(~na817_1), .IN7(~na1141_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y73     80'h00_0018_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1141_1 ( .OUT(na1141_1), .IN1(~na399_1), .IN2(1'b1), .IN3(na4293_2), .IN4(1'b1), .IN5(na2716_1), .IN6(na1029_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x42y55     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1142_4 ( .OUT(na1142_2), .IN1(~na3789_1), .IN2(~na817_1), .IN3(~na1143_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y71     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1143_1 ( .OUT(na1143_1), .IN1(na399_1), .IN2(1'b1), .IN3(~na4293_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1031_1),
                      .IN8(na2717_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x51y72     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1144_4 ( .OUT(na1144_2), .IN1(~na3792_1), .IN2(~na817_1), .IN3(~na1145_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x44y71     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1145_1 ( .OUT(na1145_1), .IN1(na399_1), .IN2(1'b1), .IN3(~na4293_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1033_1),
                      .IN8(na2718_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x39y65     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1146_1 ( .OUT(na1146_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3795_1), .IN6(~na817_1), .IN7(~na1147_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x42y67     80'h00_0018_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1147_1 ( .OUT(na1147_1), .IN1(na399_1), .IN2(1'b1), .IN3(~na4293_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1035_1),
                      .IN8(na2719_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x25y71     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1148_4 ( .OUT(na1148_2), .IN1(1'b1), .IN2(na405_2), .IN3(1'b1), .IN4(~na688_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND*/D//AND*/D      x30y79     80'h00_FE00_80_0000_0387_F858
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1149_1 ( .OUT(na1149_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3220_1), .IN6(na3231_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1149_2 ( .OUT(na1149_1), .CLK(na1739_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1149_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1149_4 ( .OUT(na1149_2_i), .IN1(na3220_1), .IN2(na3231_2), .IN3(~na1149_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1149_5 ( .OUT(na1149_2), .CLK(na1739_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1149_2_i) );
// C_MX2b/D///      x53y72     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1151_1 ( .OUT(na1151_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na3104_1), .IN7(1'b0), .IN8(na1152_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1151_2 ( .OUT(na1151_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1151_1_i) );
// C_MX2b/D///      x44y72     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1152_1 ( .OUT(na1152_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1763_2), .IN7(1'b0), .IN8(na1153_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1152_2 ( .OUT(na1152_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1152_1_i) );
// C_MX2b/D///      x44y62     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1153_1 ( .OUT(na1153_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1763_1), .IN7(1'b0), .IN8(na1154_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1153_2 ( .OUT(na1153_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1153_1_i) );
// C_MX2b/D///      x42y70     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1154_1 ( .OUT(na1154_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1765_2), .IN7(1'b0), .IN8(na1155_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1154_2 ( .OUT(na1154_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1154_1_i) );
// C_MX2b/D///      x42y68     80'h00_F600_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1155_1 ( .OUT(na1155_1_i), .IN1(~na456_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1161_1), .IN6(na1765_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1155_2 ( .OUT(na1155_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1155_1_i) );
// C_MX2b/D///      x51y73     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1156_1 ( .OUT(na1156_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1775_2), .IN7(1'b0), .IN8(na1157_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1156_2 ( .OUT(na1156_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1156_1_i) );
// C_MX2b/D///      x50y70     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1157_1 ( .OUT(na1157_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1775_1), .IN7(1'b0), .IN8(na1158_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1157_2 ( .OUT(na1157_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1157_1_i) );
// C_MX2b/D///      x48y70     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1158_1 ( .OUT(na1158_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1777_2), .IN7(1'b0), .IN8(na1159_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1158_2 ( .OUT(na1158_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1158_1_i) );
// C_MX2b/D///      x44y64     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1159_1 ( .OUT(na1159_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1777_1), .IN7(1'b0), .IN8(na1160_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1159_2 ( .OUT(na1159_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1159_1_i) );
// C_MX2b/D///      x44y54     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1160_1 ( .OUT(na1160_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4205_2), .IN5(na1161_1), .IN6(1'b0), .IN7(na3444_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1160_2 ( .OUT(na1160_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1160_1_i) );
// C_MX2b/D///      x41y53     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1161_1 ( .OUT(na1161_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4205_2), .IN5(na1162_1), .IN6(1'b0), .IN7(na3443_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1161_2 ( .OUT(na1161_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1161_1_i) );
// C_MX2b/D///      x43y53     80'h00_F600_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1162_1 ( .OUT(na1162_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4205_2), .IN5(1'b0), .IN6(na1163_1), .IN7(1'b0), .IN8(na3442_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1162_2 ( .OUT(na1162_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1162_1_i) );
// C_MX2b/D///      x45y54     80'h00_F600_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1163_1 ( .OUT(na1163_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4205_2), .IN5(1'b0), .IN6(na1164_1), .IN7(1'b0), .IN8(na3439_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1163_2 ( .OUT(na1163_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1163_1_i) );
// C_MX2b/D///      x43y54     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1164_1 ( .OUT(na1164_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4205_2), .IN5(na1165_1), .IN6(1'b0), .IN7(na3430_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1164_2 ( .OUT(na1164_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1164_1_i) );
// C_MX2b/D///      x43y55     80'h00_F600_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1165_1 ( .OUT(na1165_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4205_2), .IN5(na1603_1), .IN6(1'b0), .IN7(na3429_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1165_2 ( .OUT(na1165_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1165_1_i) );
// C_MX2b/D///      x59y78     80'h00_F600_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1166_1 ( .OUT(na1166_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4205_2), .IN5(1'b0), .IN6(na2965_1), .IN7(1'b0), .IN8(na4580_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1166_2 ( .OUT(na1166_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1166_1_i) );
// C_MX2b/D///      x56y80     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1167_1 ( .OUT(na1167_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1775_2), .IN7(1'b0), .IN8(na1168_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1167_2 ( .OUT(na1167_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1167_1_i) );
// C_MX2b/D///      x54y72     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1168_1 ( .OUT(na1168_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1767_2), .IN7(1'b0), .IN8(na1169_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1168_2 ( .OUT(na1168_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1168_1_i) );
// C_MX2b/D///      x52y72     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1169_1 ( .OUT(na1169_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1767_1), .IN7(1'b0), .IN8(na1170_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1169_2 ( .OUT(na1169_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1169_1_i) );
// C_MX2b/D///      x54y70     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1170_1 ( .OUT(na1170_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1769_2), .IN7(1'b0), .IN8(na1171_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1170_2 ( .OUT(na1170_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1170_1_i) );
// C_MX2b/D///      x50y74     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1171_1 ( .OUT(na1171_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1769_1), .IN7(1'b0), .IN8(na1172_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1171_2 ( .OUT(na1171_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1171_1_i) );
// C_MX2b/D///      x50y66     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1172_1 ( .OUT(na1172_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1771_2), .IN7(1'b0), .IN8(na1173_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1172_2 ( .OUT(na1172_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1172_1_i) );
// C_MX2b/D///      x48y64     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1173_1 ( .OUT(na1173_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1771_1), .IN7(1'b0), .IN8(na1174_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1173_2 ( .OUT(na1173_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1173_1_i) );
// C_MX2b/D///      x52y74     80'h00_F600_00_0040_0AA0_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1174_1 ( .OUT(na1174_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1773_2), .IN7(1'b0), .IN8(na1175_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1174_2 ( .OUT(na1174_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1174_1_i) );
// C_MX2b/D///      x50y76     80'h00_F600_00_0040_0AA8_00CF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1175_1 ( .OUT(na1175_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b0), .IN6(na1773_1), .IN7(1'b0), .IN8(~na1176_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1175_2 ( .OUT(na1175_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1175_1_i) );
// C_MX2b////      x54y82     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1176_1 ( .OUT(na1176_1), .IN1(1'b1), .IN2(na2965_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1156_1), .IN6(~na2965_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x31y67     80'h00_FE00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1177_1 ( .OUT(na1177_1_i), .IN1(1'b1), .IN2(~na4369_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1180_1), .IN6(na1178_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1177_2 ( .OUT(na1177_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1177_1_i) );
// C_MX2b////      x35y66     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1178_1 ( .OUT(na1178_1), .IN1(na436_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1177_1), .IN6(na1769_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x44y76     80'h00_0018_00_0000_0C88_88FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1179_1 ( .OUT(na1179_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2962_1), .IN6(na2965_2), .IN7(na2958_2),
                      .IN8(na4205_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x27y65     80'h00_FE00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1180_1 ( .OUT(na1180_1_i), .IN1(1'b1), .IN2(na4369_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1181_1), .IN8(na1182_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1180_2 ( .OUT(na1180_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1180_1_i) );
// C_MX2b////      x32y65     80'h00_0018_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1181_1 ( .OUT(na1181_1), .IN1(na436_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1180_1), .IN6(na1771_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x28y68     80'h00_FE00_00_0040_0C0A_3F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1182_1 ( .OUT(na1182_1_i), .IN1(1'b0), .IN2(na1184_1), .IN3(1'b0), .IN4(na1183_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1179_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1182_2 ( .OUT(na1182_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1182_1_i) );
// C_MX2b////      x32y66     80'h00_0018_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1183_1 ( .OUT(na1183_1), .IN1(~na436_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4475_2), .IN8(na1182_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x27y66     80'h00_FE00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1184_1 ( .OUT(na1184_1_i), .IN1(1'b1), .IN2(~na4369_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1186_1), .IN8(na1185_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1184_2 ( .OUT(na1184_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1184_1_i) );
// C_MX2b////      x34y66     80'h00_0018_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1185_1 ( .OUT(na1185_1), .IN1(~na436_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4477_2), .IN6(na1184_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x30y65     80'h00_FE00_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1186_1 ( .OUT(na1186_1_i), .IN1(na436_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1179_1), .IN5(1'b0), .IN6(1'b0), .IN7(na1186_1),
                      .IN8(na4476_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1186_2 ( .OUT(na1186_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1186_1_i) );
// C_MX4b/D///      x37y77     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1187_1 ( .OUT(na1187_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1187_1), .IN6(na30_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1187_2 ( .OUT(na1187_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1187_1_i) );
// C_MX4b/D///      x33y77     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1188_1 ( .OUT(na1188_1_i), .IN1(na1191_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1188_1), .IN6(na3943_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1188_2 ( .OUT(na1188_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1188_1_i) );
// C_MX4a////      x29y79     80'h00_0018_00_0040_0C18_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1191_1 ( .OUT(na1191_1), .IN1(1'b1), .IN2(1'b0), .IN3(1'b0), .IN4(na1296_1), .IN5(na4400_2), .IN6(1'b1), .IN7(~na287_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////D      x59y87     80'h00_FA18_00_0000_0666_3FB5
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1192_1 ( .OUT(na1192_1), .IN1(na1193_1), .IN2(1'b1), .IN3(~na3826_1), .IN4(na1388_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na1526_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1192_5 ( .OUT(na1192_2), .CLK(na1739_1), .EN(na1525_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1192_1) );
// C_AND////      x63y87     80'h00_0018_00_0000_0C88_31FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1193_1 ( .OUT(na1193_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2962_1), .IN6(~na4589_2), .IN7(1'b1), .IN8(~na1194_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x58y84     80'h00_0018_00_0000_0888_F9CC
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1194_1 ( .OUT(na1194_1), .IN1(1'b0), .IN2(~na2965_2), .IN3(1'b0), .IN4(~na1195_2), .IN5(na2962_2), .IN6(na4567_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x68y90     80'h00_0060_00_0000_0C08_FF4C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1195_4 ( .OUT(na1195_2), .IN1(1'b1), .IN2(na1196_1), .IN3(~na980_2), .IN4(na1322_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x59y92     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1196_1 ( .OUT(na1196_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na4333_2), .IN7(1'b1), .IN8(~na986_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x61y85     80'h00_0018_00_0000_0C88_CBFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1197_1 ( .OUT(na1197_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3827_1), .IN6(~na2965_2), .IN7(1'b0), .IN8(na1388_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x46y83     80'h00_F600_00_0040_0C05_4000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1198_1 ( .OUT(na1198_1_i), .IN1(na1192_1), .IN2(1'b0), .IN3(na2984_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na443_1),
                      .IN8(na450_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1198_2 ( .OUT(na1198_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1198_1_i) );
// C_ANDXOR/D//AND/D      x65y89     80'h00_FA00_80_0000_0C68_EAFA
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a1199_1 ( .OUT(na1199_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na4208_2), .IN6(1'b1), .IN7(~na2958_2),
                      .IN8(~na4627_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1199_2 ( .OUT(na1199_1), .CLK(na1739_1), .EN(na1523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1199_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1199_4 ( .OUT(na1199_2_i), .IN1(na1199_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1199_5 ( .OUT(na1199_2), .CLK(na1739_1), .EN(na1523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1199_2_i) );
// C_ORAND*/D//ORAND*/D      x41y59     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1200_1 ( .OUT(na1200_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na3098_2), .IN7(~na446_2),
                      .IN8(~na4374_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1200_2 ( .OUT(na1200_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1200_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1200_4 ( .OUT(na1200_2_i), .IN1(~na447_2), .IN2(~na3098_1), .IN3(~na446_2), .IN4(~na1202_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1200_5 ( .OUT(na1200_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1200_2_i) );
// C_ORAND*/D//ORAND*/D      x42y60     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1202_1 ( .OUT(na1202_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na3100_2), .IN7(~na446_2),
                      .IN8(~na1202_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1202_2 ( .OUT(na1202_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1202_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1202_4 ( .OUT(na1202_2_i), .IN1(~na447_2), .IN2(~na3100_1), .IN3(~na446_2), .IN4(~na4377_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1202_5 ( .OUT(na1202_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1202_2_i) );
// C_ORAND*/D//ORAND*/D      x41y62     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1204_1 ( .OUT(na1204_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na3102_2), .IN7(~na446_2),
                      .IN8(~na4378_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1204_2 ( .OUT(na1204_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1204_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1204_4 ( .OUT(na1204_2_i), .IN1(~na447_2), .IN2(~na3102_1), .IN3(~na446_2), .IN4(~na1206_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1204_5 ( .OUT(na1204_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1204_2_i) );
// C_ORAND*/D//ORAND*/D      x42y64     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1206_1 ( .OUT(na1206_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na3104_2), .IN7(~na446_2),
                      .IN8(~na1206_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1206_2 ( .OUT(na1206_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1206_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1206_4 ( .OUT(na1206_2_i), .IN1(~na447_2), .IN2(~na3104_1), .IN3(~na446_2), .IN4(~na1208_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1206_5 ( .OUT(na1206_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1206_2_i) );
// C_ORAND*/D//ORAND*/D      x38y66     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1208_1 ( .OUT(na1208_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na1763_2), .IN7(~na446_2),
                      .IN8(~na1208_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1208_2 ( .OUT(na1208_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1208_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1208_4 ( .OUT(na1208_2_i), .IN1(~na447_2), .IN2(~na1763_1), .IN3(~na446_2), .IN4(~na4381_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1208_5 ( .OUT(na1208_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1208_2_i) );
// C_ORAND*/D//ORAND*/D      x31y63     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1210_1 ( .OUT(na1210_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na1765_2), .IN7(~na446_2),
                      .IN8(~na4382_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1210_2 ( .OUT(na1210_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1210_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1210_4 ( .OUT(na1210_2_i), .IN1(~na447_2), .IN2(~na1765_1), .IN3(~na446_2), .IN4(~na1212_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1210_5 ( .OUT(na1210_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1210_2_i) );
// C_ORAND*/D//ORAND*/D      x40y64     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1212_1 ( .OUT(na1212_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na1767_2), .IN7(~na446_2),
                      .IN8(~na1212_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1212_2 ( .OUT(na1212_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1212_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1212_4 ( .OUT(na1212_2_i), .IN1(~na447_2), .IN2(~na1767_1), .IN3(~na446_2), .IN4(~na1214_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1212_5 ( .OUT(na1212_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1212_2_i) );
// C_ORAND*/D//ORAND*/D      x40y62     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1214_1 ( .OUT(na1214_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na1769_2), .IN7(~na446_2),
                      .IN8(~na1214_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1214_2 ( .OUT(na1214_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1214_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1214_4 ( .OUT(na1214_2_i), .IN1(~na447_2), .IN2(~na1769_1), .IN3(~na446_2), .IN4(~na1216_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1214_5 ( .OUT(na1214_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1214_2_i) );
// C_ORAND*/D//ORAND*/D      x38y64     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1216_1 ( .OUT(na1216_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na1771_2), .IN7(~na446_2),
                      .IN8(~na1216_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1216_2 ( .OUT(na1216_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1216_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1216_4 ( .OUT(na1216_2_i), .IN1(~na447_2), .IN2(~na1771_1), .IN3(~na446_2), .IN4(~na1218_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1216_5 ( .OUT(na1216_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1216_2_i) );
// C_ORAND*/D//ORAND*/D      x34y64     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1218_1 ( .OUT(na1218_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na1773_2), .IN7(~na446_2),
                      .IN8(~na1218_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1218_2 ( .OUT(na1218_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1218_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1218_4 ( .OUT(na1218_2_i), .IN1(~na447_2), .IN2(~na1773_1), .IN3(~na446_2), .IN4(~na1220_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1218_5 ( .OUT(na1218_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1218_2_i) );
// C_ORAND*/D//ORAND*/D      x36y64     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1220_1 ( .OUT(na1220_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na1775_2), .IN7(~na446_2),
                      .IN8(~na1220_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1220_2 ( .OUT(na1220_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1220_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1220_4 ( .OUT(na1220_2_i), .IN1(~na447_2), .IN2(~na1775_1), .IN3(~na446_2), .IN4(~na1222_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1220_5 ( .OUT(na1220_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1220_2_i) );
// C_ORAND*/D//ORAND*/D      x34y62     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1222_1 ( .OUT(na1222_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na1777_2), .IN7(~na446_2),
                      .IN8(~na1222_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1222_2 ( .OUT(na1222_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1222_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1222_4 ( .OUT(na1222_2_i), .IN1(~na447_2), .IN2(~na1777_1), .IN3(~na446_2), .IN4(~na1224_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1222_5 ( .OUT(na1222_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1222_2_i) );
// C_ORAND*/D//ORAND*/D      x36y58     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1224_1 ( .OUT(na1224_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na4602_2), .IN7(~na446_2),
                      .IN8(~na1224_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1224_2 ( .OUT(na1224_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1224_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1224_4 ( .OUT(na1224_2_i), .IN1(~na447_2), .IN2(~na4601_2), .IN3(~na446_2), .IN4(~na4392_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1224_5 ( .OUT(na1224_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1224_2_i) );
// C_ORAND*/D//ORAND*/D      x36y57     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1226_1 ( .OUT(na1226_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na4600_2), .IN7(~na446_2),
                      .IN8(~na4393_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1226_2 ( .OUT(na1226_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1226_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1226_4 ( .OUT(na1226_2_i), .IN1(~na447_2), .IN2(~na4599_2), .IN3(~na446_2), .IN4(~na1228_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1226_5 ( .OUT(na1226_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1226_2_i) );
// C_ORAND*/D//ORAND*/D      x36y56     80'h00_F600_80_0000_0387_7777
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1228_1 ( .OUT(na1228_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na4598_2), .IN7(~na446_2),
                      .IN8(~na1228_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1228_2 ( .OUT(na1228_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1228_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1228_4 ( .OUT(na1228_2_i), .IN1(~na447_2), .IN2(~na4597_2), .IN3(~na446_2), .IN4(~na4396_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1228_5 ( .OUT(na1228_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1228_2_i) );
// C_ORAND*/D//ORAND*/D      x35y53     80'h00_F600_80_0000_0387_77D7
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1230_1 ( .OUT(na1230_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na447_2), .IN6(~na4596_2), .IN7(~na446_2),
                      .IN8(~na4397_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1230_2 ( .OUT(na1230_1), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1230_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1230_4 ( .OUT(na1230_2_i), .IN1(~na447_2), .IN2(~na4595_2), .IN3(~na446_2), .IN4(na4210_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1230_5 ( .OUT(na1230_2), .CLK(na1739_1), .EN(~na1399_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1230_2_i) );
// C_///ORAND/      x66y87     80'h00_0060_00_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1232_4 ( .OUT(na1232_2), .IN1(na3895_1), .IN2(na4333_2), .IN3(~na2958_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR/D///      x32y61     80'h00_FE00_00_0000_0CEE_0D00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1233_1 ( .OUT(na1233_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na4588_2), .IN6(na1234_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1233_2 ( .OUT(na1233_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1233_1_i) );
// C_AND////      x35y70     80'h00_0018_00_0000_0888_32F2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1234_1 ( .OUT(na1234_1), .IN1(na2963_2), .IN2(~na423_1), .IN3(1'b1), .IN4(1'b1), .IN5(na3145_1), .IN6(~na423_2), .IN7(1'b1),
                      .IN8(~na1539_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x27y60     80'h00_FE00_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1235_1 ( .OUT(na1235_1_i), .IN1(1'b1), .IN2(na421_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1302_1), .IN6(na1541_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1235_2 ( .OUT(na1235_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1235_1_i) );
// C_MX2b/D///      x28y60     80'h00_FE00_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1236_1 ( .OUT(na1236_1_i), .IN1(1'b1), .IN2(na421_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1301_1), .IN6(na1541_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1236_2 ( .OUT(na1236_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1236_1_i) );
// C_///ORAND/D      x21y64     80'h00_FE00_80_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1237_4 ( .OUT(na1237_2_i), .IN1(~na3899_1), .IN2(~na421_1), .IN3(~na3898_2), .IN4(~na2971_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1237_5 ( .OUT(na1237_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1237_2_i) );
// C_ORAND/D///      x21y62     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1239_1 ( .OUT(na1239_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3902_1), .IN6(~na421_1), .IN7(~na2972_1),
                      .IN8(~na4628_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1239_2 ( .OUT(na1239_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1239_1_i) );
// C_///ORAND/D      x14y63     80'h00_FE00_80_0000_0C08_FF77
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1241_4 ( .OUT(na1241_2_i), .IN1(~na3905_1), .IN2(~na421_1), .IN3(~na3898_2), .IN4(~na4574_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1241_5 ( .OUT(na1241_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1241_2_i) );
// C_ORAND/D///      x19y59     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1243_1 ( .OUT(na1243_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3908_1), .IN6(~na421_1), .IN7(~na3898_2),
                      .IN8(~na4576_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1243_2 ( .OUT(na1243_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1243_1_i) );
// C_ORAND/D///      x21y64     80'h00_FE00_00_0000_0C88_77FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1245_1 ( .OUT(na1245_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3911_1), .IN6(~na421_1), .IN7(~na3898_2),
                      .IN8(~na4575_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1245_2 ( .OUT(na1245_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1245_1_i) );
// C_MX2b/D///      x32y50     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1247_1 ( .OUT(na1247_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4194_2), .IN5(na3912_2), .IN6(1'b0), .IN7(na3209_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1247_2 ( .OUT(na1247_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1247_1_i) );
// C_MX2b/D///      x33y50     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1248_1 ( .OUT(na1248_1_i), .IN1(1'b1), .IN2(na421_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3913_2), .IN6(na3210_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1248_2 ( .OUT(na1248_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1248_1_i) );
// C_MX2b/D///      x31y54     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1249_1 ( .OUT(na1249_1_i), .IN1(1'b1), .IN2(na421_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3914_1), .IN6(na3211_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1249_2 ( .OUT(na1249_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1249_1_i) );
// C_MX2b/D///      x33y51     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1250_1 ( .OUT(na1250_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4194_2), .IN5(na3915_1), .IN6(1'b0), .IN7(na3212_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1250_2 ( .OUT(na1250_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1250_1_i) );
// C_MX2b/D///      x33y55     80'h00_FE00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1251_1 ( .OUT(na1251_1_i), .IN1(1'b1), .IN2(~na421_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3213_1), .IN6(na3916_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1251_2 ( .OUT(na1251_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1251_1_i) );
// C_MX2b/D///      x32y53     80'h00_FE00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1252_1 ( .OUT(na1252_1_i), .IN1(1'b1), .IN2(na421_1), .IN3(1'b0), .IN4(1'b0), .IN5(na3917_2), .IN6(na3214_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1252_2 ( .OUT(na1252_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1252_1_i) );
// C_MX2b/D///      x34y58     80'h00_FE00_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1253_1 ( .OUT(na1253_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4194_2), .IN5(1'b0), .IN6(na3215_1), .IN7(1'b0), .IN8(na3918_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1253_2 ( .OUT(na1253_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1253_1_i) );
// C_ORAND*////D      x55y84     80'h00_FE18_00_0000_0788_3BB3
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1254_1 ( .OUT(na1254_1), .IN1(1'b0), .IN2(~na1260_1), .IN3(na3920_1), .IN4(~na450_1), .IN5(na1271_1), .IN6(~na1260_2), .IN7(1'b0),
                      .IN8(~na450_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1254_5 ( .OUT(na1254_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1254_1) );
// C_AND///AND/      x67y87     80'h00_0078_00_0000_0C88_415A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1255_1 ( .OUT(na1255_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2957_2), .IN6(~na4566_2), .IN7(~na2958_1),
                      .IN8(na3921_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1255_4 ( .OUT(na1255_2), .IN1(na2957_2), .IN2(1'b1), .IN3(~na2958_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ANDXOR/      x69y84     80'h00_0060_00_0000_0C06_FF5B
C_ANDXOR   #(.CPE_CFG (9'b0_1000_0000)) 
           _a1256_4 ( .OUT(na1256_2), .IN1(~na3828_1), .IN2(na1257_1), .IN3(na461_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x63y76     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1257_1 ( .OUT(na1257_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2956_1), .IN6(1'b1), .IN7(na4572_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x55y88     80'h00_0078_00_0000_0C88_8A31
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1260_1 ( .OUT(na1260_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3931_2), .IN6(1'b1), .IN7(na531_1), .IN8(na3925_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1260_4 ( .OUT(na1260_2), .IN1(~na2962_1), .IN2(~na2965_2), .IN3(1'b1), .IN4(~na4571_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x52y92     80'h00_0018_00_0000_0C88_CBFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1262_1 ( .OUT(na1262_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3927_2), .IN6(~na1263_1), .IN7(1'b0), .IN8(na532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x59y90     80'h00_0018_00_0040_0C61_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1263_1 ( .OUT(na1263_1), .IN1(na2962_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b0), .IN5(na2962_2), .IN6(1'b1), .IN7(na2961_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x55y92     80'h00_0018_00_0000_0C88_D3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1264_1 ( .OUT(na1264_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na3928_1), .IN7(~na2984_1), .IN8(na4630_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x50y89     80'h00_0018_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1269_1 ( .OUT(na1269_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1270_2), .IN6(na1528_2), .IN7(1'b0), .IN8(na532_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y85     80'h00_0060_00_0000_0C08_FF58
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1270_4 ( .OUT(na1270_2), .IN1(na507_1), .IN2(na1196_1), .IN3(~na980_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x51y79     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1271_1 ( .OUT(na1271_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na1232_2), .IN4(1'b1), .IN5(1'b0), .IN6(~na3932_1), .IN7(1'b0), .IN8(~na1605_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x65y88     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1275_1 ( .OUT(na1275_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2958_2), .IN8(na1306_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x66y84     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1276_1 ( .OUT(na1276_1), .IN1(1'b1), .IN2(na4564_2), .IN3(1'b0), .IN4(1'b0), .IN5(na3207_1), .IN6(na3208_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x34y55     80'h00_FE00_00_0040_0A50_00C0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1277_1 ( .OUT(na1277_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na4194_2), .IN5(na3938_1), .IN6(1'b0), .IN7(na3216_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1277_2 ( .OUT(na1277_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1277_1_i) );
// C_MX2b////      x29y57     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1278_1 ( .OUT(na1278_1), .IN1(1'b1), .IN2(na421_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1304_2), .IN6(na1541_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x30y58     80'h00_0018_00_0040_0A31_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1279_1 ( .OUT(na1279_1), .IN1(1'b1), .IN2(na421_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1304_1), .IN6(na1541_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x29y60     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1280_1 ( .OUT(na1280_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3899_1), .IN6(~na421_1), .IN7(~na1281_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x28y65     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1281_1 ( .OUT(na1281_1), .IN1(na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4194_2), .IN5(na1177_1), .IN6(na2966_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x25y58     80'h00_0060_00_0000_0C08_FF37
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1282_4 ( .OUT(na1282_2), .IN1(~na3902_1), .IN2(~na421_1), .IN3(1'b0), .IN4(~na1283_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x30y64     80'h00_0018_00_0040_0A30_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1283_1 ( .OUT(na1283_1), .IN1(na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4194_2), .IN5(na1180_1), .IN6(na2967_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x25y64     80'h00_0060_00_0000_0C08_FF37
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1284_4 ( .OUT(na1284_2), .IN1(~na3905_1), .IN2(~na421_1), .IN3(1'b0), .IN4(~na1285_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x28y62     80'h00_0018_00_0040_0AC0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1285_1 ( .OUT(na1285_1), .IN1(~na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4194_2), .IN5(1'b0), .IN6(1'b0), .IN7(na2968_1),
                      .IN8(na1182_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x22y62     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1286_4 ( .OUT(na1286_2), .IN1(~na3908_1), .IN2(~na421_1), .IN3(~na1287_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x26y63     80'h00_0018_00_0040_0A30_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1287_1 ( .OUT(na1287_1), .IN1(~na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4194_2), .IN5(na2969_2), .IN6(na1184_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x25y64     80'h00_0018_00_0000_0C88_37FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1288_1 ( .OUT(na1288_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3911_1), .IN6(~na421_1), .IN7(1'b0), .IN8(~na1289_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x28y58     80'h00_0018_00_0040_0AC0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1289_1 ( .OUT(na1289_1), .IN1(na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4194_2), .IN5(1'b0), .IN6(1'b0), .IN7(na1186_1),
                      .IN8(na2970_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND/D///      x33y71     80'h00_FE00_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1290_1 ( .OUT(na1290_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3940_2), .IN6(~na3939_1), .IN7(~na1149_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1290_2 ( .OUT(na1290_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1290_1_i) );
// C_MX4b/D///      x31y89     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1292_1 ( .OUT(na1292_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1292_1), .IN6(na1293_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1292_2 ( .OUT(na1292_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1292_1_i) );
// C_MX4b/D///      x29y84     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1293_1 ( .OUT(na1293_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1294_1), .IN6(na1293_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1293_2 ( .OUT(na1293_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1293_1_i) );
// C_MX4b/D///      x31y81     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1294_1 ( .OUT(na1294_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1294_1), .IN6(na1338_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1294_2 ( .OUT(na1294_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1294_1_i) );
// C_MX4b/D///      x27y79     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1295_1 ( .OUT(na1295_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1295_1), .IN6(na1298_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1295_2 ( .OUT(na1295_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1295_1_i) );
// C_ORAND/D//ORAND/D      x32y76     80'h00_FE00_80_0000_0C88_5E5E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1296_1 ( .OUT(na1296_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3307_2), .IN6(na1297_1), .IN7(~na1149_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a1296_2 ( .OUT(na1296_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1296_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1296_4 ( .OUT(na1296_2_i), .IN1(na3944_2), .IN2(na4155_2), .IN3(~na1149_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1296_5 ( .OUT(na1296_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1296_2_i) );
// C_MX4a////      x31y82     80'h00_0018_00_0040_0C29_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1297_1 ( .OUT(na1297_1), .IN1(na4631_2), .IN2(1'b1), .IN3(1'b0), .IN4(na1296_2), .IN5(1'b1), .IN6(na3943_2), .IN7(~na287_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x25y80     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1298_1 ( .OUT(na1298_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1308_1), .IN6(na1298_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1298_2 ( .OUT(na1298_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1298_1_i) );
// C_MX4b/D///      x25y67     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1301_1 ( .OUT(na1301_1_i), .IN1(1'b1), .IN2(na978_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1301_1), .IN6(na1660_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1301_2 ( .OUT(na1301_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1301_1_i) );
// C_MX4b/D///      x27y67     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1302_1 ( .OUT(na1302_1_i), .IN1(1'b1), .IN2(na978_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1302_1), .IN6(na1660_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1302_2 ( .OUT(na1302_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1302_1_i) );
// C_AND/D///      x16y62     80'h00_FE00_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1303_1 ( .OUT(na1303_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na436_1), .IN6(1'b1), .IN7(na1653_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1303_2 ( .OUT(na1303_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1303_1_i) );
// C_AND/D//AND/D      x17y63     80'h00_FE00_80_0000_0C88_C5C5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1304_1 ( .OUT(na1304_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na436_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1655_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1304_2 ( .OUT(na1304_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1304_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1304_4 ( .OUT(na1304_2_i), .IN1(~na436_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1655_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1304_5 ( .OUT(na1304_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1304_2_i) );
// C_///AND/D      x26y51     80'h00_FE00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1305_4 ( .OUT(na1305_2_i), .IN1(na888_2), .IN2(1'b1), .IN3(1'b1), .IN4(na3426_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1305_5 ( .OUT(na1305_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1305_2_i) );
// C_AND/D//ORAND*/D      x66y90     80'h00_FE00_80_0000_0C87_5AB3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1306_1 ( .OUT(na1306_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1637_1), .IN6(1'b1), .IN7(~na443_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1306_2 ( .OUT(na1306_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1306_1_i) );
C_ORAND    #(.CPE_CFG (9'b1_1000_0000)) 
           _a1306_4 ( .OUT(na1306_2_i), .IN1(1'b0), .IN2(~na4402_2), .IN3(na2958_2), .IN4(~na4457_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1306_5 ( .OUT(na1306_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1306_2_i) );
// C_AND/D//AND/D      x65y92     80'h00_FE00_80_0000_0C88_5C5C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1307_1 ( .OUT(na1307_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1635_2), .IN7(~na443_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1307_2 ( .OUT(na1307_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1307_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1307_4 ( .OUT(na1307_2_i), .IN1(1'b1), .IN2(na1635_1), .IN3(~na443_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1307_5 ( .OUT(na1307_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1307_2_i) );
// C_MX4b/D///      x27y81     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1308_1 ( .OUT(na1308_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1308_1), .IN6(na1312_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1308_2 ( .OUT(na1308_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1308_1_i) );
// C_MX4b/D///      x32y81     80'h00_FE00_00_0040_0AC8_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1309_1 ( .OUT(na1309_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1309_1),
                      .IN8(~na1310_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1309_2 ( .OUT(na1309_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1309_1_i) );
// C_MX2b////      x48y88     80'h00_0018_00_0040_0ACC_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1310_1 ( .OUT(na1310_1), .IN1(na457_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1269_1), .IN8(~na1311_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x50y86     80'h00_0060_00_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1311_4 ( .OUT(na1311_2), .IN1(1'b1), .IN2(1'b1), .IN3(na531_1), .IN4(na3925_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x29y82     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1312_1 ( .OUT(na1312_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na4403_2), .IN6(na1312_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1312_2 ( .OUT(na1312_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1312_1_i) );
// C_MX4b/D///      x30y84     80'h00_FE00_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1313_1 ( .OUT(na1313_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1336_1),
                      .IN8(na1313_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1313_2 ( .OUT(na1313_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1313_1_i) );
// C_///ORAND/D      x59y65     80'h00_FE00_80_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1314_4 ( .OUT(na1314_2_i), .IN1(na3948_1), .IN2(na1315_2), .IN3(~na1149_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a1314_5 ( .OUT(na1314_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1314_2_i) );
// C_///ORAND/      x31y68     80'h00_0060_00_0000_0C08_FFEC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1315_4 ( .OUT(na1315_2), .IN1(1'b0), .IN2(na137_2), .IN3(na3950_2), .IN4(na420_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x14y73     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1316_1 ( .OUT(na1316_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na318_1), .IN8(~na420_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x25y84     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1317_1 ( .OUT(na1317_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na727_1), .IN6(na1317_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1317_2 ( .OUT(na1317_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1317_1_i) );
// C_MX4b/D///      x25y82     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1318_1 ( .OUT(na1318_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na692_1), .IN6(na1318_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1318_2 ( .OUT(na1318_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1318_1_i) );
// C_MX4b/D///      x21y73     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1319_1 ( .OUT(na1319_1_i), .IN1(1'b1), .IN2(na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na1319_1), .IN6(na640_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1319_2 ( .OUT(na1319_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1319_1_i) );
// C_MX4b/D///      x19y74     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1320_1 ( .OUT(na1320_1_i), .IN1(1'b1), .IN2(~na424_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na4254_2), .IN6(na1320_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1320_2 ( .OUT(na1320_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1320_1_i) );
// C_MX4b/D///      x51y88     80'h00_FE00_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1321_1 ( .OUT(na1321_1_i), .IN1(na456_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4404_2),
                      .IN8(na1322_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1321_2 ( .OUT(na1321_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1321_1_i) );
// C_MX4b/D///      x54y88     80'h00_FE00_00_0040_0AC3_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1322_1 ( .OUT(na1322_1_i), .IN1(~na456_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na4214_2),
                      .IN8(na1322_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1322_2 ( .OUT(na1322_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1322_1_i) );
// C_MX4b/D///      x26y90     80'h00_FE00_00_0040_0AC0_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1323_1 ( .OUT(na1323_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4405_2),
                      .IN8(na1323_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1323_2 ( .OUT(na1323_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1323_1_i) );
// C_MX4b/D///      x25y88     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1324_1 ( .OUT(na1324_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1327_1), .IN6(na1324_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1324_2 ( .OUT(na1324_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1324_1_i) );
// C_MX4b/D///      x43y88     80'h00_FE00_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1325_1 ( .OUT(na1325_1_i), .IN1(na430_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4406_2),
                      .IN8(na1683_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1325_2 ( .OUT(na1325_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1325_1_i) );
// C_MX4b/D///      x44y89     80'h00_FE00_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1326_1 ( .OUT(na1326_1_i), .IN1(na430_2), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1326_1),
                      .IN8(na1683_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1326_2 ( .OUT(na1326_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1326_1_i) );
// C_MX4b/D///      x27y85     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1327_1 ( .OUT(na1327_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1327_1), .IN6(na1328_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1327_2 ( .OUT(na1327_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1327_1_i) );
// C_MX4b/D///      x27y86     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1328_1 ( .OUT(na1328_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1329_1), .IN6(na1328_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1328_2 ( .OUT(na1328_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1328_1_i) );
// C_MX4b/D///      x29y89     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1329_1 ( .OUT(na1329_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1329_1), .IN6(na1331_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1329_2 ( .OUT(na1329_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1329_1_i) );
// C_AND/D//AND/D      x48y86     80'h00_FE00_80_0000_0C88_A5A5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1330_1 ( .OUT(na1330_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na218_1), .IN6(1'b1), .IN7(na1680_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1330_2 ( .OUT(na1330_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1330_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1330_4 ( .OUT(na1330_2_i), .IN1(~na218_1), .IN2(1'b1), .IN3(na1680_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1330_5 ( .OUT(na1330_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1330_2_i) );
// C_MX4b/D///      x31y88     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1331_1 ( .OUT(na1331_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na4410_2), .IN6(na1352_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1331_2 ( .OUT(na1331_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1331_1_i) );
// C_MX4b/D///      x28y90     80'h00_FE00_00_0040_0AC4_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1332_1 ( .OUT(na1332_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1333_1),
                      .IN8(na1332_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1332_2 ( .OUT(na1332_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1332_1_i) );
// C_MX2b////      x32y87     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1333_1 ( .OUT(na1333_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1341_2), .IN5(1'b0), .IN6(~na1334_2), .IN7(1'b0), .IN8(~na1127_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x35y84     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1334_4 ( .OUT(na1334_2), .IN1(na3809_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1337_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x27y89     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1335_1 ( .OUT(na1335_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1335_1), .IN6(na1376_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1335_2 ( .OUT(na1335_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1335_1_i) );
// C_MX4b/D///      x28y83     80'h00_FE00_00_0040_0AC0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1336_1 ( .OUT(na1336_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1336_1),
                      .IN8(na1323_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1336_2 ( .OUT(na1336_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1336_1_i) );
// C_ORAND*/D///      x34y84     80'h00_FE00_00_0000_0788_5FB5
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1337_1 ( .OUT(na1337_1_i), .IN1(~na220_1), .IN2(1'b0), .IN3(na1517_2), .IN4(~na1337_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na1149_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1337_2 ( .OUT(na1337_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1337_1_i) );
// C_MX4b/D///      x29y80     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1338_1 ( .OUT(na1338_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1295_1), .IN6(na1338_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1338_2 ( .OUT(na1338_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1338_1_i) );
// C_MX4b/D///      x45y75     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1339_1 ( .OUT(na1339_1_i), .IN1(na31_2), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1339_1), .IN6(na44_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1339_2 ( .OUT(na1339_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1339_1_i) );
// C_MX4b/D///      x34y85     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1340_1 ( .OUT(na1340_1_i), .IN1(1'b1), .IN2(na232_1), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1340_1),
                      .IN8(na1347_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1340_2 ( .OUT(na1340_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1340_1_i) );
// C_///ORAND/D      x38y86     80'h00_FE00_80_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1341_4 ( .OUT(na1341_2_i), .IN1(na3954_1), .IN2(na1342_1), .IN3(~na1149_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1341_5 ( .OUT(na1341_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1341_2_i) );
// C_MX4a////      x37y88     80'h00_0018_00_0040_0C82_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1342_1 ( .OUT(na1342_1), .IN1(1'b0), .IN2(na3955_2), .IN3(1'b0), .IN4(1'b1), .IN5(na1345_1), .IN6(1'b1), .IN7(na2713_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x45y91     80'h00_0018_00_0040_0C55_1000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1343_1 ( .OUT(na1343_1), .IN1(~na1037_1), .IN2(1'b0), .IN3(~na1344_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na4545_2),
                      .IN8(~na2707_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x42y85     80'h00_0060_00_0000_0C08_FF6C
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1344_4 ( .OUT(na1344_2), .IN1(1'b0), .IN2(~na1509_2), .IN3(~na1038_1), .IN4(na993_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x33y85     80'h00_0018_00_0000_0C88_84FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1345_1 ( .OUT(na1345_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2712_2), .IN6(na232_2), .IN7(na2713_1),
                      .IN8(na1347_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x34y89     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1346_1 ( .OUT(na1346_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na232_2), .IN7(1'b1), .IN8(na1347_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1346_2 ( .OUT(na1346_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1346_1_i) );
// C_MX4b/D///      x30y92     80'h00_FE00_00_0040_0AC4_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1347_1 ( .OUT(na1347_1_i), .IN1(1'b1), .IN2(~na4412_2), .IN3(~na4141_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1349_1),
                      .IN8(na1347_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1347_2 ( .OUT(na1347_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1347_1_i) );
// C_AND///AND/      x34y91     80'h00_0078_00_0000_0C88_C15A
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1349_1 ( .OUT(na1349_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1118_2), .IN6(~na225_2), .IN7(1'b1), .IN8(na229_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1349_4 ( .OUT(na1349_2), .IN1(na222_1), .IN2(1'b1), .IN3(~na1340_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x22y82     80'h00_F600_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1350_4 ( .OUT(na1350_2_i), .IN1(na411_1), .IN2(na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1350_5 ( .OUT(na1350_2), .CLK(na1739_1), .EN(~na1418_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1350_2_i) );
// C_///ORAND/D      x26y83     80'h00_FE00_80_0000_0C08_FFE3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1351_4 ( .OUT(na1351_2_i), .IN1(1'b0), .IN2(~na288_2), .IN3(na1351_2), .IN4(na3958_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1351_5 ( .OUT(na1351_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1351_2_i) );
// C_MX4b/D///      x29y86     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1352_1 ( .OUT(na1352_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1335_1), .IN6(na1352_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1352_2 ( .OUT(na1352_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1352_1_i) );
// C_MX4b/D///      x15y54     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1353_1 ( .OUT(na1353_1_i), .IN1(~na212_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1716_2), .IN6(na1353_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1353_2 ( .OUT(na1353_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1353_1_i) );
// C_AND/D///      x45y81     80'h00_FE00_00_0000_0888_5122
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1354_1 ( .OUT(na1354_1_i), .IN1(na820_1), .IN2(~na285_1), .IN3(na83_2), .IN4(~na3230_2), .IN5(~na1354_1), .IN6(~na285_2),
                      .IN7(~na1149_2), .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1354_2 ( .OUT(na1354_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1354_1_i) );
// C_MX4b/D///      x19y79     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1355_1 ( .OUT(na1355_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na1355_1), .IN6(na4117_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1355_2 ( .OUT(na1355_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1355_1_i) );
// C_MX4b/D///      x19y80     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1356_1 ( .OUT(na1356_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na163_1), .IN6(na1356_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1356_2 ( .OUT(na1356_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1356_1_i) );
// C_MX4b/D///      x21y79     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1357_1 ( .OUT(na1357_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na1357_1), .IN6(na1356_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1357_2 ( .OUT(na1357_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1357_1_i) );
// C_MX2b/D///      x30y54     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1358_1 ( .OUT(na1358_1_i), .IN1(~na888_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3443_2), .IN8(na1359_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1358_2 ( .OUT(na1358_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1358_1_i) );
// C_MX2b/D///      x24y48     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1359_1 ( .OUT(na1359_1_i), .IN1(na888_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1360_1), .IN8(na3442_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1359_2 ( .OUT(na1359_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1359_1_i) );
// C_MX2b/D///      x24y45     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1360_1 ( .OUT(na1360_1_i), .IN1(na888_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1361_1), .IN8(na3439_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1360_2 ( .OUT(na1360_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1360_1_i) );
// C_MX2b/D///      x24y47     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1361_1 ( .OUT(na1361_1_i), .IN1(~na888_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3430_1), .IN8(na1362_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1361_2 ( .OUT(na1361_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1361_1_i) );
// C_MX2b/D///      x26y48     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1362_1 ( .OUT(na1362_1_i), .IN1(~na888_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3429_2), .IN8(na1363_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1362_2 ( .OUT(na1362_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1362_1_i) );
// C_MX2b/D///      x28y50     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1363_1 ( .OUT(na1363_1_i), .IN1(na888_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1305_2), .IN8(na3427_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1363_2 ( .OUT(na1363_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1363_1_i) );
// C_MX4b/D///      x19y81     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1364_1 ( .OUT(na1364_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na1364_1), .IN6(na158_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1364_2 ( .OUT(na1364_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1364_1_i) );
// C_MX4b/D///      x18y78     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1365_1 ( .OUT(na1365_1_i), .IN1(1'b1), .IN2(~na120_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na134_1),
                      .IN8(na1365_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1365_2 ( .OUT(na1365_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1365_1_i) );
// C_MX4b/D///      x19y69     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1366_1 ( .OUT(na1366_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na1366_1), .IN6(na130_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1366_2 ( .OUT(na1366_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1366_1_i) );
// C_MX4b/D///      x19y67     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1367_1 ( .OUT(na1367_1_i), .IN1(1'b1), .IN2(na120_2), .IN3(na1149_2), .IN4(1'b1), .IN5(na1367_1), .IN6(na4415_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1367_2 ( .OUT(na1367_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1367_1_i) );
// C_MX4b/D///      x29y91     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1368_1 ( .OUT(na1368_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1368_1), .IN6(na1377_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1368_2 ( .OUT(na1368_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1368_1_i) );
// C_MX4b/D///      x20y63     80'h00_FE00_00_0040_0AC3_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1369_1 ( .OUT(na1369_1_i), .IN1(1'b1), .IN2(na1487_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1369_1),
                      .IN8(na4100_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1369_2 ( .OUT(na1369_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1369_1_i) );
// C_///ORAND/D      x27y69     80'h00_FE00_80_0000_0C08_FF5E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1370_4 ( .OUT(na1370_2_i), .IN1(na1371_1), .IN2(na3960_2), .IN3(~na1149_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1370_5 ( .OUT(na1370_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1370_2_i) );
// C_MX4a////      x21y61     80'h00_0018_00_0040_0C41_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1371_1 ( .OUT(na1371_1), .IN1(na3961_2), .IN2(1'b0), .IN3(1'b1), .IN4(1'b0), .IN5(~na1374_2), .IN6(1'b1), .IN7(na4529_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x23y65     80'h00_0018_00_0040_0C33_0100
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1372_1 ( .OUT(na1372_1), .IN1(~na877_1), .IN2(~na1373_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na4521_2), .IN6(~na2474_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x19y52     80'h00_0060_00_0000_0C08_FF6C
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1373_4 ( .OUT(na1373_2), .IN1(1'b0), .IN2(~na1487_1), .IN3(~na4298_2), .IN4(na864_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x15y61     80'h00_0060_00_0000_0C08_FF82
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1374_4 ( .OUT(na1374_2), .IN1(na4163_2), .IN2(~na2478_1), .IN3(na2481_2), .IN4(na214_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x15y53     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1375_4 ( .OUT(na1375_2_i), .IN1(1'b1), .IN2(na299_1), .IN3(1'b1), .IN4(na214_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1375_5 ( .OUT(na1375_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1375_2_i) );
// C_MX4b/D///      x29y88     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1376_1 ( .OUT(na1376_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1368_1), .IN6(na1376_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1376_2 ( .OUT(na1376_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1376_1_i) );
// C_MX4b/D///      x31y86     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1377_1 ( .OUT(na1377_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na4417_2), .IN6(na1381_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1377_2 ( .OUT(na1377_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1377_1_i) );
// C_MX4b/D///      x25y87     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1378_1 ( .OUT(na1378_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1378_1), .IN6(na1379_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1378_2 ( .OUT(na1378_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1378_1_i) );
// C_MX4b/D///      x23y86     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1379_1 ( .OUT(na1379_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1397_1), .IN6(na1379_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1379_2 ( .OUT(na1379_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1379_1_i) );
// C_MX4b/D///      x27y82     80'h00_FE00_00_0040_0A30_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1381_1 ( .OUT(na1381_1_i), .IN1(~na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1378_1), .IN6(na1381_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1381_2 ( .OUT(na1381_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1381_1_i) );
// C_///ORAND/D      x47y56     80'h00_FE00_80_0000_0C08_FFAE
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1383_4 ( .OUT(na1383_2_i), .IN1(na335_2), .IN2(na1383_2), .IN3(na3964_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1383_5 ( .OUT(na1383_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1383_2_i) );
// C_OR/D//OR/D      x16y86     80'h00_FE00_80_0000_0CEE_AEBC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1385_1 ( .OUT(na1385_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1618_2), .IN6(na288_2), .IN7(na287_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1385_2 ( .OUT(na1385_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1385_1_i) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a1385_4 ( .OUT(na1385_2_i), .IN1(1'b0), .IN2(na288_2), .IN3(na287_2), .IN4(~na1385_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1385_5 ( .OUT(na1385_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1385_2_i) );
// C_MX4b/D///      x43y62     80'h00_FE00_00_0040_0AC0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1386_1 ( .OUT(na1386_1_i), .IN1(1'b1), .IN2(~na1383_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1730_1),
                      .IN8(na4418_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1386_2 ( .OUT(na1386_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1386_1_i) );
// C_MX4b/D///      x45y63     80'h00_FE00_00_0040_0AC0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1387_1 ( .OUT(na1387_1_i), .IN1(1'b1), .IN2(na1383_2), .IN3(~na1149_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na4419_2),
                      .IN8(na1728_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1387_2 ( .OUT(na1387_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1387_1_i) );
// C_MX2b/D///      x56y74     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1388_1 ( .OUT(na1388_1_i), .IN1(~na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3444_1), .IN8(na1389_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1388_2 ( .OUT(na1388_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1388_1_i) );
// C_MX2b/D///      x34y52     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1389_1 ( .OUT(na1389_1_i), .IN1(~na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3443_2), .IN8(na1390_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1389_2 ( .OUT(na1389_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1389_1_i) );
// C_MX2b/D///      x32y54     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1390_1 ( .OUT(na1390_1_i), .IN1(na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1391_1), .IN8(na3442_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1390_2 ( .OUT(na1390_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1390_1_i) );
// C_MX2b/D///      x26y47     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1391_1 ( .OUT(na1391_1_i), .IN1(na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1392_1), .IN8(na3439_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1391_2 ( .OUT(na1391_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1391_1_i) );
// C_MX2b/D///      x26y49     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1392_1 ( .OUT(na1392_1_i), .IN1(~na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3430_1), .IN8(na1393_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1392_2 ( .OUT(na1392_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1392_1_i) );
// C_MX2b/D///      x28y52     80'h00_FE00_00_0040_0AC0_00F5
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1393_1 ( .OUT(na1393_1_i), .IN1(~na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na3429_2), .IN8(na1394_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1393_2 ( .OUT(na1393_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1393_1_i) );
// C_MX2b/D///      x32y52     80'h00_FE00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1394_1 ( .OUT(na1394_1_i), .IN1(na888_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na887_2), .IN8(na3427_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1394_2 ( .OUT(na1394_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1394_1_i) );
// C_MX4b/D///      x29y75     80'h00_FE00_00_0040_0A30_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1395_1 ( .OUT(na1395_1_i), .IN1(1'b1), .IN2(na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1395_1), .IN6(na4168_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1395_2 ( .OUT(na1395_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1395_1_i) );
// C_MX4b/D///      x27y74     80'h00_FE00_00_0040_0A30_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1396_1 ( .OUT(na1396_1_i), .IN1(1'b1), .IN2(~na33_1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1395_1), .IN6(na1396_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1396_2 ( .OUT(na1396_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1396_1_i) );
// C_MX4b/D///      x25y85     80'h00_FE00_00_0040_0A30_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1397_1 ( .OUT(na1397_1_i), .IN1(na220_1), .IN2(1'b1), .IN3(na1149_2), .IN4(1'b1), .IN5(na1397_1), .IN6(na361_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1397_2 ( .OUT(na1397_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1397_1_i) );
// C_ORAND////      x38y74     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1398_1 ( .OUT(na1398_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4399_2), .IN6(~na4401_2), .IN7(~na287_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x40y63     80'h00_0018_00_0000_0C88_ADFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1399_1 ( .OUT(na1399_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na456_1), .IN6(na4584_2), .IN7(na446_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x47y66     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1400_1 ( .OUT(na1400_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na436_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na4205_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x60y78     80'h00_0060_00_0000_0C08_FFDC
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1401_4 ( .OUT(na1401_2), .IN1(1'b0), .IN2(na223_2), .IN3(~na4140_2), .IN4(na3285_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x49y75     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1402_4 ( .OUT(na1402_2), .IN1(~na218_1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x22y46     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1403_1 ( .OUT(na1403_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na121_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na4442_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x43y48     80'h00_0018_00_0000_0C88_BAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1404_1 ( .OUT(na1404_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na301_1), .IN6(1'b0), .IN7(na4587_2), .IN8(~na4442_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x58y57     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1405_4 ( .OUT(na1405_2), .IN1(1'b1), .IN2(~na4424_2), .IN3(1'b1), .IN4(~na54_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x69y49     80'h00_0060_00_0000_0C08_FFCB
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1406_4 ( .OUT(na1406_2), .IN1(na4585_2), .IN2(~na4424_2), .IN3(1'b0), .IN4(na4091_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x66y42     80'h00_0018_00_0000_0C88_CDFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1407_1 ( .OUT(na1407_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1465_2), .IN6(na4586_2), .IN7(1'b0), .IN8(na336_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y45     80'h00_0018_00_0000_0C88_35FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1408_1 ( .OUT(na1408_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na275_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na4432_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y52     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1409_1 ( .OUT(na1409_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4467_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1544_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x61y47     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1410_1 ( .OUT(na1410_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4467_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1544_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x62y48     80'h00_0018_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1411_1 ( .OUT(na1411_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4467_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1544_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y40     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1412_1 ( .OUT(na1412_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4464_2), .IN6(~na1542_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x61y40     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1413_1 ( .OUT(na1413_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4464_2), .IN6(na1542_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y36     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1414_4 ( .OUT(na1414_2), .IN1(na4464_2), .IN2(na1542_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x36y46     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1415_4 ( .OUT(na1415_2), .IN1(na4468_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1545_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x39y46     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1416_1 ( .OUT(na1416_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4468_2), .IN6(1'b1), .IN7(1'b1), .IN8(na1545_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x36y48     80'h00_0060_00_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1417_4 ( .OUT(na1417_2), .IN1(na4468_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1545_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x29y87     80'h00_0060_00_0000_0C08_FF73
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1418_4 ( .OUT(na1418_2), .IN1(1'b0), .IN2(~na288_2), .IN3(~na287_2), .IN4(~na1296_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x57y70     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1419_4 ( .OUT(na1419_2), .IN1(na4466_2), .IN2(~na1543_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x51y75     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1420_1 ( .OUT(na1420_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4466_2), .IN6(na1543_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x51y76     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1421_1 ( .OUT(na1421_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4466_2), .IN6(na1543_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x39y59     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1422_1 ( .OUT(na1422_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1541_1), .IN7(1'b1), .IN8(na4462_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x39y59     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1423_4 ( .OUT(na1423_2), .IN1(1'b1), .IN2(na1541_1), .IN3(1'b1), .IN4(~na4462_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x32y57     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1424_4 ( .OUT(na1424_2), .IN1(1'b1), .IN2(na1541_1), .IN3(1'b1), .IN4(na4462_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x68y64     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1425_4 ( .OUT(na1425_2), .IN1(1'b1), .IN2(~na2350_2), .IN3(1'b1), .IN4(~na519_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x69y45     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1426_4 ( .OUT(na1426_2), .IN1(~na704_2), .IN2(~na2246_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x39y55     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1427_4 ( .OUT(na1427_2), .IN1(1'b1), .IN2(~na881_2), .IN3(1'b1), .IN4(~na2497_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x53y92     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1428_1 ( .OUT(na1428_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1044_2), .IN7(1'b1), .IN8(~na2730_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y81     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1429_4 ( .OUT(na1429_2), .IN1(~na1192_2), .IN2(~na2981_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x36y55     80'h00_0018_00_0000_0C88_D3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1431_1 ( .OUT(na1431_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na4424_2), .IN7(~na4093_2), .IN8(na1090_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x61y64     80'h00_FE00_00_0000_0C88_34FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1432_1 ( .OUT(na1432_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na3975_1), .IN6(na4075_2), .IN7(1'b1), .IN8(~na1434_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1432_2 ( .OUT(na1432_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1432_1_i) );
// C_MX4b////      x66y70     80'h00_0018_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1434_1 ( .OUT(na1434_1), .IN1(na4489_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1990_1), .IN5(na4490_2), .IN6(~na1993_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x66y79     80'h00_0018_00_0000_0888_FDAC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1435_1 ( .OUT(na1435_1), .IN1(1'b0), .IN2(na523_1), .IN3(na115_1), .IN4(1'b0), .IN5(~na360_2), .IN6(na103_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x67y79     80'h00_0060_00_0000_0C08_FF84
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1436_4 ( .OUT(na1436_2), .IN1(~na360_2), .IN2(na57_1), .IN3(na115_1), .IN4(na4222_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x70y75     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1437_1 ( .OUT(na1437_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na522_2), .IN6(1'b1), .IN7(na115_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x69y76     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1438_1 ( .OUT(na1438_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3977_1), .IN7(na115_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1438_2 ( .OUT(na1438_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1438_1_i) );
// C_AND/D///      x66y81     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1439_1 ( .OUT(na1439_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na31_2), .IN6(na3978_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1439_2 ( .OUT(na1439_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1439_1_i) );
// C_///AND/D      x64y88     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1440_4 ( .OUT(na1440_2_i), .IN1(na31_2), .IN2(na3979_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1440_5 ( .OUT(na1440_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1440_2_i) );
// C_///AND/D      x67y62     80'h00_FA00_80_0000_0C08_FFC8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1441_4 ( .OUT(na1441_2_i), .IN1(na535_1), .IN2(na1986_2), .IN3(1'b1), .IN4(na1984_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1441_5 ( .OUT(na1441_2), .CLK(na1739_1), .EN(na115_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1441_2_i) );
// C_AND*/D//ORAND/D      x58y64     80'h00_FE00_80_0000_0388_3C5E
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1443_1 ( .OUT(na1443_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4424_2), .IN7(1'b1), .IN8(~na1088_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1443_2 ( .OUT(na1443_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1443_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1443_4 ( .OUT(na1443_2_i), .IN1(na90_1), .IN2(na4424_2), .IN3(~na38_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1443_5 ( .OUT(na1443_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1443_2_i) );
// C_AND/D///      x66y67     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1444_1 ( .OUT(na1444_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4424_2), .IN7(na511_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1444_2 ( .OUT(na1444_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1444_1_i) );
// C_MX4a////D      x69y77     80'h00_FA18_00_0040_0C49_A300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1445_1 ( .OUT(na1445_1), .IN1(na4426_2), .IN2(1'b0), .IN3(1'b1), .IN4(na1446_2), .IN5(1'b1), .IN6(~na512_1), .IN7(na4221_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1445_5 ( .OUT(na1445_2), .CLK(na1739_1), .EN(na1435_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1445_1) );
// C_///AND/D      x70y76     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1446_4 ( .OUT(na1446_2_i), .IN1(na1445_1), .IN2(na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1446_5 ( .OUT(na1446_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1446_2_i) );
// C_AND/D///      x66y65     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1447_1 ( .OUT(na1447_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3981_1), .IN6(na4424_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1447_2 ( .OUT(na1447_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1447_1_i) );
// C_ORAND////      x70y65     80'h00_0018_00_0000_0C88_E3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1448_1 ( .OUT(na1448_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na1986_1), .IN7(na3983_1), .IN8(na519_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x69y66     80'h00_0060_00_0000_0C08_FFB3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1449_4 ( .OUT(na1449_2), .IN1(1'b0), .IN2(~na1986_1), .IN3(na4519_2), .IN4(~na519_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x69y67     80'h00_0060_00_0000_0C08_FFB3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1450_4 ( .OUT(na1450_2), .IN1(1'b0), .IN2(~na1986_1), .IN3(na3983_1), .IN4(~na519_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x57y58     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1451_1 ( .OUT(na1451_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4223_2), .IN7(1'b1), .IN8(na1411_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1451_2 ( .OUT(na1451_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1451_1_i) );
// C_///ORAND/      x23y56     80'h00_0060_00_0000_0C08_FFB5
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1453_4 ( .OUT(na1453_2), .IN1(~na1465_2), .IN2(1'b0), .IN3(na4179_2), .IN4(~na340_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x52y55     80'h00_FE00_80_0000_0C08_FF34
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1454_4 ( .OUT(na1454_2_i), .IN1(~na1456_1), .IN2(na33_1), .IN3(1'b1), .IN4(~na3988_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1454_5 ( .OUT(na1454_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1454_2_i) );
// C_MX4b////      x53y61     80'h00_0018_00_0040_0A51_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1456_1 ( .OUT(na1456_1), .IN1(1'b1), .IN2(na2228_2), .IN3(1'b1), .IN4(~na4511_2), .IN5(~na2229_1), .IN6(1'b0), .IN7(na4506_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x49y61     80'h00_0018_00_0000_0888_FBAA
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1457_1 ( .OUT(na1457_1), .IN1(na333_1), .IN2(1'b0), .IN3(na262_1), .IN4(1'b0), .IN5(na329_1), .IN6(~na295_1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x53y63     80'h00_0060_00_0000_0C08_FF28
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1458_4 ( .OUT(na1458_2), .IN1(na333_1), .IN2(na330_1), .IN3(na262_1), .IN4(~na4159_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x55y64     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1459_4 ( .OUT(na1459_2), .IN1(na707_1), .IN2(na4173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x64y60     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1460_4 ( .OUT(na1460_2_i), .IN1(na3990_1), .IN2(na4173_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1460_5 ( .OUT(na1460_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1460_2_i) );
// C_AND/D///      x60y72     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1461_1 ( .OUT(na1461_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3991_1), .IN7(1'b1), .IN8(na4076_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1461_2 ( .OUT(na1461_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1461_1_i) );
// C_///AND/D      x54y75     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1462_4 ( .OUT(na1462_2_i), .IN1(na3992_1), .IN2(na33_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1462_5 ( .OUT(na1462_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1462_2_i) );
// C_AND/D///      x65y47     80'h00_FA00_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1463_1 ( .OUT(na1463_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4265_2), .IN6(1'b1), .IN7(na2223_2), .IN8(na2221_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1463_2 ( .OUT(na1463_1), .CLK(na1739_1), .EN(na333_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1463_1_i) );
// C_AND*/D//ORAND/D      x55y55     80'h00_FE00_80_0000_0388_5A3E
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1465_1 ( .OUT(na1465_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1465_2), .IN6(1'b1), .IN7(~na356_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1465_2 ( .OUT(na1465_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1465_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1465_4 ( .OUT(na1465_2_i), .IN1(na1465_2), .IN2(na4174_2), .IN3(1'b0), .IN4(~na4160_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1465_5 ( .OUT(na1465_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1465_2_i) );
// C_AND/D///      x63y52     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1466_1 ( .OUT(na1466_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1465_2), .IN6(na352_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1466_2 ( .OUT(na1466_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1466_1_i) );
// C_MX4a////D      x56y63     80'h00_FA18_00_0040_0C86_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1467_1 ( .OUT(na1467_1), .IN1(1'b0), .IN2(na4435_2), .IN3(na1468_1), .IN4(1'b1), .IN5(na707_1), .IN6(1'b1), .IN7(na353_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1467_5 ( .OUT(na1467_2), .CLK(na1739_1), .EN(na1457_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1467_1) );
// C_AND/D///      x54y59     80'h00_FE00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1468_1 ( .OUT(na1468_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1465_2), .IN6(1'b1), .IN7(na1467_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1468_2 ( .OUT(na1468_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1468_1_i) );
// C_AND/D///      x62y49     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1469_1 ( .OUT(na1469_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1465_2), .IN6(na3994_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1469_2 ( .OUT(na1469_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1469_1_i) );
// C_ORAND////      x69y46     80'h00_0018_00_0000_0C88_5EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1470_1 ( .OUT(na1470_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3996_2), .IN6(na2246_2), .IN7(~na2223_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x68y47     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1471_4 ( .OUT(na1471_2), .IN1(na704_2), .IN2(~na2246_2), .IN3(~na2223_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x70y48     80'h00_0018_00_0000_0C88_5BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1472_1 ( .OUT(na1472_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3996_2), .IN6(~na2246_2), .IN7(~na2223_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x51y41     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1473_4 ( .OUT(na1473_2_i), .IN1(1'b1), .IN2(na1414_2), .IN3(na636_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1473_5 ( .OUT(na1473_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1473_2_i) );
// C_ORAND////      x18y42     80'h00_0018_00_0000_0C88_3BFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1475_1 ( .OUT(na1475_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1375_2), .IN6(~na4165_2), .IN7(1'b0), .IN8(~na4442_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x13y56     80'h00_FE00_80_0000_0C08_FF34
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1476_4 ( .OUT(na1476_2_i), .IN1(~na1478_1), .IN2(na120_2), .IN3(1'b1), .IN4(~na4001_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1476_5 ( .OUT(na1476_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1476_2_i) );
// C_MX4b////      x17y55     80'h00_0018_00_0040_0AC4_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1478_1 ( .OUT(na1478_1), .IN1(1'b1), .IN2(~na2478_2), .IN3(~na4526_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na2481_2),
                      .IN8(na4532_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x15y55     80'h00_0018_00_0000_0888_BFAC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1479_1 ( .OUT(na1479_1), .IN1(1'b0), .IN2(na299_1), .IN3(na189_2), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na1369_1), .IN8(~na214_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x22y64     80'h00_0018_00_0000_0C88_84FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1480_1 ( .OUT(na1480_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4131_2), .IN6(na299_1), .IN7(na189_2), .IN8(na110_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x21y55     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1481_4 ( .OUT(na1481_2), .IN1(1'b1), .IN2(na299_1), .IN3(1'b1), .IN4(na884_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x15y62     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1482_4 ( .OUT(na1482_2_i), .IN1(1'b1), .IN2(na299_1), .IN3(na4003_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1482_5 ( .OUT(na1482_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1482_2_i) );
// C_///AND/D      x13y67     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1483_4 ( .OUT(na1483_2_i), .IN1(1'b1), .IN2(na4004_1), .IN3(na4104_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1483_5 ( .OUT(na1483_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1483_2_i) );
// C_///AND/D      x15y71     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1484_4 ( .OUT(na1484_2_i), .IN1(1'b1), .IN2(na4005_1), .IN3(na4104_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1484_5 ( .OUT(na1484_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1484_2_i) );
// C_AND/D///      x28y51     80'h00_FA00_00_0000_0C88_C8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1485_1 ( .OUT(na1485_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2472_1), .IN6(na2474_2), .IN7(1'b1), .IN8(na864_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1485_2 ( .OUT(na1485_1), .CLK(na1739_1), .EN(na299_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1485_1_i) );
// C_AND*/D//ORAND/D      x25y54     80'h00_FE00_80_0000_0388_C3E3
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1487_1 ( .OUT(na1487_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1373_2), .IN7(1'b1), .IN8(na4442_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1487_2 ( .OUT(na1487_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1487_1_i) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1487_4 ( .OUT(na1487_2_i), .IN1(1'b0), .IN2(~na4132_2), .IN3(na1567_1), .IN4(na4442_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1487_5 ( .OUT(na1487_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1487_2_i) );
// C_AND/D///      x23y59     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1488_1 ( .OUT(na1488_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na877_1), .IN6(1'b1), .IN7(1'b1), .IN8(na4442_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1488_2 ( .OUT(na1488_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1488_1_i) );
// C_MX4a////D      x18y50     80'h00_FA18_00_0040_0C29_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1489_1 ( .OUT(na1489_1), .IN1(na1490_2), .IN2(1'b1), .IN3(1'b0), .IN4(na4445_2), .IN5(1'b1), .IN6(na878_1), .IN7(1'b1), .IN8(~na884_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1489_5 ( .OUT(na1489_2), .CLK(na1739_1), .EN(na1479_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1489_1) );
// C_///AND/D      x15y49     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1490_4 ( .OUT(na1490_2_i), .IN1(1'b1), .IN2(na4441_2), .IN3(1'b1), .IN4(na1489_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1490_5 ( .OUT(na1490_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1490_2_i) );
// C_AND/D///      x24y55     80'h00_FE00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1491_1 ( .OUT(na1491_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1487_2), .IN7(1'b1), .IN8(na4007_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1491_2 ( .OUT(na1491_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1491_1_i) );
// C_ORAND////      x35y50     80'h00_0018_00_0000_0C88_E3FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1492_1 ( .OUT(na1492_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(~na2474_1), .IN7(na4009_1), .IN8(na2497_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x36y55     80'h00_0060_00_0000_0C08_FFB3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1493_4 ( .OUT(na1493_2), .IN1(1'b0), .IN2(~na2474_1), .IN3(na4302_2), .IN4(~na2497_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x42y56     80'h00_0060_00_0000_0C08_FFB3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1494_4 ( .OUT(na1494_2), .IN1(1'b0), .IN2(~na2474_1), .IN3(na4009_1), .IN4(~na2497_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x26y54     80'h00_FE00_80_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1495_4 ( .OUT(na1495_2_i), .IN1(1'b1), .IN2(na194_1), .IN3(1'b1), .IN4(na1417_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1495_5 ( .OUT(na1495_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1495_2_i) );
// C_///ORAND/      x25y89     80'h00_0060_00_0000_0C08_FFB3
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1497_4 ( .OUT(na1497_2), .IN1(1'b0), .IN2(~na232_1), .IN3(na1346_1), .IN4(~na4139_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x35y81     80'h00_FE00_00_0000_0C88_1AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1498_1 ( .OUT(na1498_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na220_1), .IN6(1'b1), .IN7(~na1500_1), .IN8(~na4014_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1498_2 ( .OUT(na1498_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1498_1_i) );
// C_MX4b////      x36y83     80'h00_0018_00_0040_0A54_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1500_1 ( .OUT(na1500_1), .IN1(na2712_2), .IN2(1'b1), .IN3(na2713_2), .IN4(1'b1), .IN5(na2712_1), .IN6(1'b0), .IN7(~na2713_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x28y91     80'h00_0018_00_0000_0888_DFCC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1501_1 ( .OUT(na1501_1), .IN1(1'b0), .IN2(na1048_1), .IN3(1'b0), .IN4(na1347_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na432_2),
                      .IN8(na239_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x39y92     80'h00_0018_00_0000_0C88_84FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1502_1 ( .OUT(na1502_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4198_2), .IN6(na1048_1), .IN7(na238_1),
                      .IN8(na1347_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x39y92     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1503_4 ( .OUT(na1503_2), .IN1(1'b1), .IN2(na1047_1), .IN3(1'b1), .IN4(na1347_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x41y90     80'h00_FE00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1504_4 ( .OUT(na1504_2_i), .IN1(na4411_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4016_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1504_5 ( .OUT(na1504_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1504_2_i) );
// C_///AND/D      x31y90     80'h00_FE00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1505_4 ( .OUT(na1505_2_i), .IN1(na4017_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4137_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1505_5 ( .OUT(na1505_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1505_2_i) );
// C_AND/D///      x25y90     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1506_1 ( .OUT(na1506_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4018_1), .IN6(1'b1), .IN7(1'b1), .IN8(na4137_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1506_2 ( .OUT(na1506_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1506_1_i) );
// C_AND/D///      x36y81     80'h00_FA00_00_0000_0C88_8AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1507_1 ( .OUT(na1507_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4547_2), .IN6(1'b1), .IN7(na2705_2), .IN8(na993_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1507_2 ( .OUT(na1507_1), .CLK(na1739_1), .EN(na1347_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1507_1_i) );
// C_///AND*/D      x39y84     80'h00_FE00_80_0000_0C07_FF5C
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1509_4 ( .OUT(na1509_2_i), .IN1(1'b1), .IN2(na232_1), .IN3(~na1344_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1509_5 ( .OUT(na1509_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1509_2_i) );
// C_AND/D///      x37y87     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1510_1 ( .OUT(na1510_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1037_1), .IN6(na232_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1510_2 ( .OUT(na1510_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1510_1_i) );
// C_MX4a////D      x36y89     80'h00_FA18_00_0040_0C29_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1511_1 ( .OUT(na1511_1), .IN1(na4451_2), .IN2(1'b1), .IN3(1'b0), .IN4(na1512_1), .IN5(1'b1), .IN6(na1047_1), .IN7(~na1038_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1511_5 ( .OUT(na1511_2), .CLK(na1739_1), .EN(na1501_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1511_1) );
// C_AND/D///      x36y90     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1512_1 ( .OUT(na1512_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na232_1), .IN7(na1511_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1512_2 ( .OUT(na1512_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1512_1_i) );
// C_AND/D///      x35y84     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1513_1 ( .OUT(na1513_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4020_1), .IN6(na232_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1513_2 ( .OUT(na1513_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1513_1_i) );
// C_///ORAND/      x55y91     80'h00_0060_00_0000_0C08_FF3E
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1514_4 ( .OUT(na1514_2), .IN1(na4558_2), .IN2(na4022_2), .IN3(1'b0), .IN4(~na2707_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x54y92     80'h00_0060_00_0000_0C08_FF3D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1515_4 ( .OUT(na1515_2), .IN1(~na4558_2), .IN2(na1044_2), .IN3(1'b0), .IN4(~na2707_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x56y89     80'h00_0060_00_0000_0C08_FF3D
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1516_4 ( .OUT(na1516_2), .IN1(~na4558_2), .IN2(na4022_2), .IN3(1'b0), .IN4(~na2707_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x52y81     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1517_4 ( .OUT(na1517_2_i), .IN1(1'b1), .IN2(na1421_1), .IN3(na4293_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1517_5 ( .OUT(na1517_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1517_2_i) );
// C_ORAND////      x18y75     80'h00_0018_00_0000_0C88_D5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1519_1 ( .OUT(na1519_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na456_1), .IN6(1'b0), .IN7(~na449_2), .IN8(na4212_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/D      x37y71     80'h00_FE00_80_0000_0C08_FF43
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1520_4 ( .OUT(na1520_2_i), .IN1(1'b1), .IN2(~na4027_1), .IN3(~na1522_1), .IN4(na4195_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1520_5 ( .OUT(na1520_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1520_2_i) );
// C_MX4b////      x54y83     80'h00_0018_00_0040_0A32_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1522_1 ( .OUT(na1522_1), .IN1(na2962_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4568_2), .IN5(na2963_2), .IN6(~na2965_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x61y91     80'h00_0018_00_0000_0888_DFAC
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1523_1 ( .OUT(na1523_1), .IN1(1'b0), .IN2(na1196_1), .IN3(na443_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(~na980_2), .IN8(na1322_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x62y88     80'h00_0060_00_0000_0C08_FF48
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1524_4 ( .OUT(na1524_2), .IN1(na4371_2), .IN2(na1321_1), .IN3(~na980_2), .IN4(na4201_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x62y88     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1525_1 ( .OUT(na1525_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na443_1), .IN8(na1195_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x64y88     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1526_1 ( .OUT(na1526_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na4029_1), .IN7(na443_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1526_2 ( .OUT(na1526_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1526_1_i) );
// C_///AND/D      x52y91     80'h00_FE00_80_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1527_4 ( .OUT(na1527_2_i), .IN1(na4030_1), .IN2(na424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1527_5 ( .OUT(na1527_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1527_2_i) );
// C_///AND/D      x43y90     80'h00_FE00_80_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1528_4 ( .OUT(na1528_2_i), .IN1(1'b1), .IN2(na424_2), .IN3(na4031_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1528_5 ( .OUT(na1528_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1528_2_i) );
// C_///AND/D      x62y78     80'h00_FA00_80_0000_0C08_FF8A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1529_4 ( .OUT(na1529_2_i), .IN1(na2956_1), .IN2(1'b1), .IN3(na2958_2), .IN4(na1388_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1529_5 ( .OUT(na1529_2), .CLK(na1739_1), .EN(na443_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1529_2_i) );
// C_///AND*/D      x63y79     80'h00_FE00_80_0000_0C07_FF5A
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1531_4 ( .OUT(na1531_2_i), .IN1(na456_1), .IN2(1'b1), .IN3(~na467_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1531_5 ( .OUT(na1531_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1531_2_i) );
// C_AND/D///      x61y81     80'h00_FE00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1532_1 ( .OUT(na1532_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na460_1), .IN6(1'b1), .IN7(1'b1), .IN8(na4205_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1532_2 ( .OUT(na1532_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1532_1_i) );
// C_MX4a////D      x67y85     80'h00_FA18_00_0040_0C86_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1533_1 ( .OUT(na1533_1), .IN1(1'b0), .IN2(na4458_2), .IN3(na1534_2), .IN4(1'b1), .IN5(1'b1), .IN6(na4209_2), .IN7(1'b1),
                      .IN8(na1195_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1533_5 ( .OUT(na1533_2), .CLK(na1739_1), .EN(na1523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1533_1) );
// C_///AND/D      x70y87     80'h00_FE00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1534_4 ( .OUT(na1534_2_i), .IN1(na1533_1), .IN2(1'b1), .IN3(1'b1), .IN4(na4205_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1534_5 ( .OUT(na1534_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1534_2_i) );
// C_AND/D///      x63y79     80'h00_FE00_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1535_1 ( .OUT(na1535_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na456_1), .IN6(na4033_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1535_2 ( .OUT(na1535_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1535_1_i) );
// C_ORAND////      x59y86     80'h00_0018_00_0000_0C88_5EFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1536_1 ( .OUT(na1536_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4035_2), .IN6(na2981_1), .IN7(~na2958_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x66y81     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1537_4 ( .OUT(na1537_2), .IN1(na1192_2), .IN2(~na2981_1), .IN3(~na2958_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x64y84     80'h00_0060_00_0000_0C08_FF5B
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1538_4 ( .OUT(na1538_2), .IN1(na4035_2), .IN2(~na2981_1), .IN3(~na2958_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x30y66     80'h00_FE00_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1539_1 ( .OUT(na1539_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na421_1), .IN7(na1424_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1539_2 ( .OUT(na1539_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1539_1_i) );
// C_///AND/      x13y71     80'h00_0060_00_0000_0C08_FF1F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1540_4 ( .OUT(na1540_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na990_1), .IN4(~na1350_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR/D//AND/D      x31y62     80'h00_FA00_80_0000_0C68_CCF3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1541_1 ( .OUT(na1541_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1541_1), .IN7(1'b0), .IN8(na4462_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1541_2 ( .OUT(na1541_1), .CLK(na1739_1), .EN(na421_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1541_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1541_4 ( .OUT(na1541_2_i), .IN1(1'b1), .IN2(~na1541_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1541_5 ( .OUT(na1541_2), .CLK(na1739_1), .EN(na421_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1541_2_i) );
// C_XOR/D//AND/D      x69y36     80'h00_FA00_80_0000_0C68_06F3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1542_1 ( .OUT(na1542_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4464_2), .IN6(na1542_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1542_2 ( .OUT(na1542_1), .CLK(na1739_1), .EN(na636_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1542_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1542_4 ( .OUT(na1542_2_i), .IN1(1'b1), .IN2(~na1542_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1542_5 ( .OUT(na1542_2), .CLK(na1739_1), .EN(na636_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1542_2_i) );
// C_XOR/D//AND/D      x55y78     80'h00_FA00_80_0000_0C68_06F3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1543_1 ( .OUT(na1543_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4466_2), .IN6(na1543_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1543_2 ( .OUT(na1543_1), .CLK(na1739_1), .EN(na817_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1543_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1543_4 ( .OUT(na1543_2_i), .IN1(1'b1), .IN2(~na1543_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1543_5 ( .OUT(na1543_2), .CLK(na1739_1), .EN(na817_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1543_2_i) );
// C_XOR/D//AND/D      x68y46     80'h00_FA00_80_0000_0C68_CA3F
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1544_1 ( .OUT(na1544_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4467_2), .IN6(1'b0), .IN7(1'b0), .IN8(na1544_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1544_2 ( .OUT(na1544_1), .CLK(na1739_1), .EN(na526_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1544_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1544_4 ( .OUT(na1544_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1544_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1544_5 ( .OUT(na1544_2), .CLK(na1739_1), .EN(na526_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1544_2_i) );
// C_XOR/D//AND/D      x40y48     80'h00_FA00_80_0000_0C68_CA3F
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1545_1 ( .OUT(na1545_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4468_2), .IN6(1'b0), .IN7(1'b0), .IN8(na1545_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1545_2 ( .OUT(na1545_1), .CLK(na1739_1), .EN(na194_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1545_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1545_4 ( .OUT(na1545_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1545_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1545_5 ( .OUT(na1545_2), .CLK(na1739_1), .EN(na194_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1545_2_i) );
// C_OR////      x23y91     80'h00_0018_00_0000_0EEE_7577
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1564_1 ( .OUT(na1564_1), .IN1(~na4045_2), .IN2(~na225_2), .IN3(~na1340_1), .IN4(~na3268_1), .IN5(~na4045_1), .IN6(1'b0),
                      .IN7(~na4046_1), .IN8(~na3268_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND*////D      x20y53     80'h00_FE18_00_0000_0788_CB3B
C_ORAND    #(.CPE_CFG (9'b1_0000_0000)) 
           _a1567_1 ( .OUT(na1567_1), .IN1(na301_1), .IN2(~na957_2), .IN3(1'b0), .IN4(~na200_1), .IN5(na307_1), .IN6(~na4416_2), .IN7(1'b0),
                      .IN8(na1608_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1567_5 ( .OUT(na1567_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1567_1) );
// C_OR////      x44y53     80'h00_0018_00_0000_0EEE_5777
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1570_1 ( .OUT(na1570_1), .IN1(~na3296_1), .IN2(~na4053_2), .IN3(~na4054_2), .IN4(~na340_2), .IN5(~na3296_2), .IN6(~na4053_1),
                      .IN7(~na332_1), .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x64y89     80'h00_0018_00_0000_0EEE_7757
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1574_1 ( .OUT(na1574_1), .IN1(~na3322_1), .IN2(~na4058_2), .IN3(~na449_2), .IN4(1'b0), .IN5(~na3322_2), .IN6(~na4058_1),
                      .IN7(~na4059_2), .IN8(~na518_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x64y72     80'h00_0018_00_0040_0C98_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1576_1 ( .OUT(na1576_1), .IN1(1'b1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1990_1), .IN5(1'b1), .IN6(~na1989_2), .IN7(1'b1), .IN8(na1990_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x64y67     80'h00_0018_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1577_1 ( .OUT(na1577_1), .IN1(~na4489_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1576_1), .IN5(na486_1), .IN6(na1993_1), .IN7(na4491_2),
                      .IN8(na4213_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x66y63     80'h00_0018_00_0040_0C0C_F400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1578_1 ( .OUT(na1578_1), .IN1(1'b0), .IN2(1'b0), .IN3(na1577_1), .IN4(na485_1), .IN5(~na4489_2), .IN6(na1993_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x49y53     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1579_1 ( .OUT(na1579_1_i), .IN1(1'b1), .IN2(~na4424_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1578_1), .IN8(na3712_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1579_2 ( .OUT(na1579_1), .CLK(na1739_1), .EN(~na1405_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1579_1_i) );
// C_MX4a////      x70y59     80'h00_0018_00_0040_0C43_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1580_1 ( .OUT(na1580_1), .IN1(na567_1), .IN2(na559_1), .IN3(1'b1), .IN4(1'b0), .IN5(1'b1), .IN6(~na2350_2), .IN7(1'b1), .IN8(~na519_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////D      x70y64     80'h00_F618_00_0040_0A58_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1581_1 ( .OUT(na1581_1), .IN1(1'b1), .IN2(na4220_2), .IN3(na1580_1), .IN4(1'b1), .IN5(na543_1), .IN6(1'b0), .IN7(na551_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1581_5 ( .OUT(na1581_2), .CLK(na1739_1), .EN(~na575_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1581_1) );
// C_MX4a////      x62y60     80'h00_0018_00_0040_0C62_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1582_1 ( .OUT(na1582_1), .IN1(1'b0), .IN2(~na2228_2), .IN3(1'b1), .IN4(1'b0), .IN5(na2229_2), .IN6(1'b1), .IN7(na2226_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y59     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1583_1 ( .OUT(na1583_1), .IN1(na2229_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1582_1), .IN5(na4512_2), .IN6(na664_1), .IN7(na4257_2),
                      .IN8(na2230_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x53y58     80'h00_0018_00_0040_0C03_0400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1584_1 ( .OUT(na1584_1), .IN1(na1583_1), .IN2(na663_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2229_2), .IN6(na4509_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x48y44     80'h00_F600_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1585_1 ( .OUT(na1585_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4432_2), .IN5(1'b0), .IN6(na1584_1), .IN7(1'b0), .IN8(na3720_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1585_2 ( .OUT(na1585_1), .CLK(na1739_1), .EN(~na1408_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1585_1_i) );
// C_MX4a////      x72y44     80'h00_0018_00_0040_0C25_5300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1586_1 ( .OUT(na1586_1), .IN1(na752_1), .IN2(1'b1), .IN3(na744_1), .IN4(1'b0), .IN5(1'b1), .IN6(~na2246_2), .IN7(~na4261_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////D      x71y44     80'h00_F618_00_0040_0A58_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1587_1 ( .OUT(na1587_1), .IN1(1'b1), .IN2(na2246_2), .IN3(1'b1), .IN4(na1586_1), .IN5(na4267_2), .IN6(1'b0), .IN7(na736_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1587_5 ( .OUT(na1587_2), .CLK(na1739_1), .EN(~na761_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1587_1) );
// C_MX4a////      x14y53     80'h00_0018_00_0040_0C62_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1588_1 ( .OUT(na1588_1), .IN1(1'b0), .IN2(~na2478_1), .IN3(1'b1), .IN4(1'b0), .IN5(1'b1), .IN6(na2478_2), .IN7(1'b1), .IN8(na4525_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x17y49     80'h00_0018_00_0040_0AF0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1589_1 ( .OUT(na1589_1), .IN1(1'b1), .IN2(~na2478_2), .IN3(na1588_1), .IN4(1'b1), .IN5(na843_1), .IN6(na4533_2), .IN7(na2481_1),
                      .IN8(na4295_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x21y46     80'h00_0018_00_0040_0C03_0200
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1590_1 ( .OUT(na1590_1), .IN1(na1589_1), .IN2(na842_1), .IN3(1'b0), .IN4(1'b0), .IN5(na4534_2), .IN6(~na2478_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x22y42     80'h00_F600_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1591_1 ( .OUT(na1591_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na4442_2), .IN5(1'b0), .IN6(na1590_1), .IN7(1'b0), .IN8(na3526_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1591_2 ( .OUT(na1591_1), .CLK(na1739_1), .EN(~na1403_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1591_1_i) );
// C_MX4a////      x41y51     80'h00_0018_00_0040_0C83_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1592_1 ( .OUT(na1592_1), .IN1(na908_1), .IN2(na916_1), .IN3(1'b0), .IN4(1'b1), .IN5(1'b1), .IN6(na881_2), .IN7(1'b1), .IN8(~na2497_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////D      x39y52     80'h00_F618_00_0040_0A38_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1593_1 ( .OUT(na1593_1), .IN1(na1592_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2497_1), .IN5(na4304_2), .IN6(na900_1), .IN7(1'b0),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1593_5 ( .OUT(na1593_2), .CLK(na1739_1), .EN(~na924_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1593_1) );
// C_MX4a////      x40y83     80'h00_0018_00_0040_0C91_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1594_1 ( .OUT(na1594_1), .IN1(~na2712_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b1), .IN5(1'b1), .IN6(~na4553_2), .IN7(1'b1), .IN8(na2710_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x41y79     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1595_1 ( .OUT(na1595_1), .IN1(1'b1), .IN2(na4553_2), .IN3(na1594_1), .IN4(1'b1), .IN5(na2714_1), .IN6(na1016_1), .IN7(na4336_2),
                      .IN8(na4554_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x38y77     80'h00_0018_00_0040_0C05_4000
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1596_1 ( .OUT(na1596_1), .IN1(na1595_1), .IN2(1'b0), .IN3(na1015_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na2713_2),
                      .IN8(na4552_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x36y68     80'h00_F600_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1597_1 ( .OUT(na1597_1_i), .IN1(1'b1), .IN2(~na232_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1596_1), .IN8(na3414_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1597_2 ( .OUT(na1597_1), .CLK(na1739_1), .EN(~na1402_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1597_1_i) );
// C_MX4a////      x57y85     80'h00_0018_00_0040_0C43_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1598_1 ( .OUT(na1598_1), .IN1(na1076_1), .IN2(na4350_2), .IN3(1'b1), .IN4(1'b0), .IN5(1'b1), .IN6(~na1044_2), .IN7(1'b1),
                      .IN8(~na2730_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////D      x54y85     80'h00_F618_00_0040_0A34_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1599_1 ( .OUT(na1599_1), .IN1(~na1598_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2730_2), .IN5(na1060_1), .IN6(na1052_1), .IN7(1'b1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1599_5 ( .OUT(na1599_2), .CLK(na1739_1), .EN(~na1084_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1599_1) );
// C_MX4a////      x58y89     80'h00_0018_00_0040_0C91_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1600_1 ( .OUT(na1600_1), .IN1(~na2962_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b1), .IN5(~na2962_2), .IN6(1'b1), .IN7(na2961_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y83     80'h00_0018_00_0040_0AF0_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1601_1 ( .OUT(na1601_1), .IN1(~na2962_2), .IN2(1'b1), .IN3(na1600_1), .IN4(1'b1), .IN5(na4368_2), .IN6(na2965_1), .IN7(na4573_2),
                      .IN8(na1167_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x56y79     80'h00_0018_00_0040_0C03_0400
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1602_1 ( .OUT(na1602_1), .IN1(na1601_1), .IN2(na1166_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2962_2), .IN6(na2965_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a/D///      x43y59     80'h00_F600_00_0040_0C0C_F500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1603_1 ( .OUT(na1603_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1602_1), .IN4(na3427_1), .IN5(~na456_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1603_2 ( .OUT(na1603_1), .CLK(na1739_1), .EN(~na1400_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1603_1_i) );
// C_MX4a////      x52y73     80'h00_0018_00_0040_0C1C_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1604_1 ( .OUT(na1604_1), .IN1(1'b1), .IN2(1'b0), .IN3(na4391_2), .IN4(na1216_1), .IN5(~na1192_2), .IN6(1'b1), .IN7(na4577_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////D      x54y78     80'h00_F618_00_0040_0AA4_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1605_1 ( .OUT(na1605_1), .IN1(1'b1), .IN2(~na2981_1), .IN3(na1604_1), .IN4(1'b1), .IN5(1'b0), .IN6(na4373_2), .IN7(1'b1),
                      .IN8(na1208_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1605_5 ( .OUT(na1605_2), .CLK(na1739_1), .EN(~na1232_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1605_1) );
// C_OR////      x14y54     80'h00_0018_00_0000_0EEE_7775
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a1608_1 ( .OUT(na1608_1), .IN1(~na4063_1), .IN2(1'b0), .IN3(~na4050_1), .IN4(~na303_2), .IN5(~na4063_2), .IN6(~na4064_1),
                      .IN7(~na4050_2), .IN8(~na124_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x14y62     80'h00_0078_00_0020_0C66_530C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1610_1 ( .OUT(na1610_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na2_2), .IN7(~na318_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1612_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1610_4 ( .OUT(na1610_2), .COUTY1(na1610_4), .IN1(1'b1), .IN2(na2_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na2_2), .IN7(~na318_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na1612_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x14y61     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1612_2 ( .OUT(na1612_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1612_6 ( .COUTY1(na1612_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1612_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x14y63     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a1613_1 ( .OUT(na1613_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1610_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x13y59     80'h00_0078_00_0020_0C66_A3C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1614_1 ( .OUT(na1614_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na405_2), .IN7(na317_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1616_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1614_4 ( .OUT(na1614_2), .COUTY1(na1614_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na26_1), .IN5(1'b1), .IN6(~na405_2),
                      .IN7(na317_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1616_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x13y58     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1616_2 ( .OUT(na1616_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1616_6 ( .COUTY1(na1616_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1616_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x13y60     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a1617_1 ( .OUT(na1617_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1614_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x15y83     80'h00_0078_00_0020_0C66_CCCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1618_1 ( .OUT(na1618_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na288_1), .IN7(1'b1), .IN8(na1385_2),
                      .CINX(1'b0), .CINY1(na1627_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1618_4 ( .OUT(na1618_2), .COUTY1(na1618_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1385_1), .IN5(1'b1), .IN6(na288_1),
                      .IN7(1'b1), .IN8(na1385_2), .CINX(1'b0), .CINY1(na1627_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x15y84     80'h00_0078_00_0020_0C66_AFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1620_1 ( .OUT(na1620_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na287_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1618_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1620_4 ( .OUT(na1620_2), .COUTY1(na1620_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na289_1), .IN5(1'b1), .IN6(1'b1), .IN7(na287_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na1618_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x15y85     80'h00_0078_00_0020_0C66_CFCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1622_1 ( .OUT(na1622_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na292_2),
                      .CINX(1'b0), .CINY1(na1620_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1622_4 ( .OUT(na1622_2), .COUTY1(na1622_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na292_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na292_2), .CINX(1'b0), .CINY1(na1620_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x15y86     80'h00_0078_00_0020_0C66_FCAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1624_1 ( .OUT(na1624_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na293_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1622_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1624_4 ( .OUT(na1624_2), .COUTY1(na1624_4), .IN1(1'b1), .IN2(1'b1), .IN3(na294_2), .IN4(1'b1), .IN5(1'b1), .IN6(na293_2),
                      .IN7(1'b1), .IN8(1'b1), .CINX(1'b0), .CINY1(na1622_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x15y87     80'h00_0018_00_0010_0666_00FC
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1626_1 ( .OUT(na1626_1), .IN1(1'b1), .IN2(na288_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1624_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x15y82     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1627_2 ( .OUT(na1627_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1627_6 ( .COUTY1(na1627_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1627_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x60y76     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1628_1 ( .OUT(na1628_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4095_2), .IN6(1'b1), .IN7(1'b1), .IN8(na104_1),
                      .CINX(1'b0), .CINY1(na1632_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1628_4 ( .OUT(na1628_2), .COUTY1(na1628_4), .IN1(na109_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4095_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na104_1), .CINX(1'b0), .CINY1(na1632_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x60y77     80'h00_0078_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1630_1 ( .OUT(na1630_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na428_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1628_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1630_4 ( .OUT(na1630_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na108_1), .IN5(1'b1), .IN6(na428_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1628_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x60y75     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1632_2 ( .OUT(na1632_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1632_6 ( .COUTY1(na1632_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1632_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x67y89     80'h00_0078_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1633_1 ( .OUT(na1633_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na825_1), .IN7(1'b1), .IN8(na826_2),
                      .CINX(1'b0), .CINY1(na1638_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1633_4 ( .OUT(na1633_2), .COUTY1(na1633_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na826_1), .IN5(1'b1), .IN6(na825_1),
                      .IN7(1'b1), .IN8(na826_2), .CINX(1'b0), .CINY1(na1638_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x67y90     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1635_1 ( .OUT(na1635_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1307_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1633_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1635_4 ( .OUT(na1635_2), .COUTY1(na1635_4), .IN1(1'b1), .IN2(na1307_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1307_2),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1633_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x67y91     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1637_1 ( .OUT(na1637_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1306_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1635_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x67y88     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1638_2 ( .OUT(na1638_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1638_6 ( .COUTY1(na1638_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1638_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x63y48     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1639_1 ( .OUT(na1639_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na88_2), .IN7(na87_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1648_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1639_4 ( .OUT(na1639_2), .COUTY1(na1639_4), .IN1(1'b1), .IN2(na88_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na88_2), .IN7(na87_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(na1648_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x63y49     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1641_1 ( .OUT(na1641_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na89_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1639_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1641_4 ( .OUT(na1641_2), .IN1(1'b1), .IN2(na89_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na89_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1639_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x64y81     80'h00_0078_00_0020_0C66_AA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1643_1 ( .OUT(na1643_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na360_2), .IN6(1'b1), .IN7(na246_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1652_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1643_4 ( .OUT(na1643_2), .COUTY1(na1643_4), .IN1(na360_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na360_2), .IN6(1'b1),
                      .IN7(na246_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na1652_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x64y82     80'h00_0018_00_0010_0666_00A0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1645_1 ( .OUT(na1645_1), .IN1(1'b0), .IN2(1'b0), .IN3(na38_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1643_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x52y80     80'h00_0078_00_0020_0C66_CACC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1646_1 ( .OUT(na1646_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1192_2), .IN6(1'b1), .IN7(1'b1), .IN8(na986_2),
                      .CINX(1'b0), .CINY1(na1657_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1646_4 ( .OUT(na1646_2), .COUTY1(na1646_4), .IN1(1'b1), .IN2(na2981_1), .IN3(1'b1), .IN4(na986_1), .IN5(na1192_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na986_2), .CINX(1'b0), .CINY1(na1657_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x63y47     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1648_2 ( .OUT(na1648_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1648_6 ( .COUTY1(na1648_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1648_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x56y90     80'h00_0078_00_0020_0C66_ACC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1649_1 ( .OUT(na1649_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na510_1), .IN7(na980_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1664_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1649_4 ( .OUT(na1649_2), .COUTY1(na1649_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na986_2), .IN5(1'b1), .IN6(na510_1),
                      .IN7(na980_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1664_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x56y91     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1651_1 ( .OUT(na1651_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na986_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1649_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x64y80     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1652_2 ( .OUT(na1652_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1652_6 ( .COUTY1(na1652_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1652_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x14y57     80'h00_0078_00_0020_0C66_CC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1653_1 ( .OUT(na1653_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na927_2), .IN7(1'b1), .IN8(na1303_1),
                      .CINX(1'b0), .CINY1(na1665_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1653_4 ( .OUT(na1653_2), .COUTY1(na1653_4), .IN1(1'b1), .IN2(na927_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na927_2),
                      .IN7(1'b1), .IN8(na1303_1), .CINX(1'b0), .CINY1(na1665_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x14y58     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1655_1 ( .OUT(na1655_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1304_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1653_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1655_4 ( .OUT(na1655_2), .IN1(na1304_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1304_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1653_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x52y79     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1657_2 ( .OUT(na1657_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1657_6 ( .COUTY1(na1657_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1657_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x31y71     80'h00_0078_00_0020_0C66_CA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1658_1 ( .OUT(na1658_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4331_2), .IN6(1'b1), .IN7(1'b1), .IN8(na926_1),
                      .CINX(1'b0), .CINY1(na1673_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1658_4 ( .OUT(na1658_2), .COUTY1(na1658_4), .IN1(1'b1), .IN2(na929_1), .IN3(1'b0), .IN4(1'b0), .IN5(na4331_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na926_1), .CINX(1'b0), .CINY1(na1673_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x31y72     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1660_1 ( .OUT(na1660_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1302_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1658_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1660_4 ( .OUT(na1660_2), .IN1(na1301_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1302_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1658_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x67y69     80'h00_0078_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1662_1 ( .OUT(na1662_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na360_1), .IN6(1'b1), .IN7(na4519_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1677_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1662_4 ( .OUT(na1662_2), .COUTY1(na1662_4), .IN1(na4077_2), .IN2(1'b1), .IN3(1'b1), .IN4(na519_2), .IN5(na360_1), .IN6(1'b1),
                      .IN7(na4519_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1677_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x56y89     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1664_2 ( .OUT(na1664_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1664_6 ( .COUTY1(na1664_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1664_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x14y56     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1665_2 ( .OUT(na1665_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1665_6 ( .COUTY1(na1665_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1665_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x17y89     80'h00_0078_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1666_1 ( .OUT(na1666_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na387_2), .IN7(na388_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1682_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1666_4 ( .OUT(na1666_2), .COUTY1(na1666_4), .IN1(1'b0), .IN2(1'b0), .IN3(na388_1), .IN4(1'b1), .IN5(1'b1), .IN6(na387_2),
                      .IN7(na388_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1682_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x17y90     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1668_1 ( .OUT(na1668_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na390_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1666_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1668_4 ( .OUT(na1668_2), .COUTY1(na1668_4), .IN1(na390_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na390_2), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1666_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x17y91     80'h00_0018_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1670_1 ( .OUT(na1670_1), .IN1(1'b1), .IN2(na391_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1668_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x46y89     80'h00_0078_00_0020_0C66_CACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1671_1 ( .OUT(na1671_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na434_2), .IN6(1'b1), .IN7(1'b1), .IN8(na4340_2),
                      .CINX(1'b0), .CINY1(na1687_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1671_4 ( .OUT(na1671_2), .COUTY1(na1671_4), .IN1(na434_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2730_2), .IN5(na434_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na4340_2), .CINX(1'b0), .CINY1(na1687_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x31y70     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1673_2 ( .OUT(na1673_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1673_6 ( .COUTY1(na1673_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1673_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x30y88     80'h00_0078_00_0020_0C66_AA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1674_1 ( .OUT(na1674_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4145_2), .IN6(1'b1), .IN7(na432_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1693_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1674_4 ( .OUT(na1674_2), .COUTY1(na1674_4), .IN1(na434_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na4145_2), .IN6(1'b1),
                      .IN7(na432_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1693_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x30y89     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1676_1 ( .OUT(na1676_1), .IN1(na434_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1674_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x67y68     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1677_2 ( .OUT(na1677_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1677_6 ( .COUTY1(na1677_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1677_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x44y84     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1678_1 ( .OUT(na1678_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na403_2), .IN7(na402_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1701_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1678_4 ( .OUT(na1678_2), .COUTY1(na1678_4), .IN1(1'b1), .IN2(na403_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na403_2),
                      .IN7(na402_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1701_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x44y85     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1680_1 ( .OUT(na1680_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1330_2),
                      .CINX(1'b0), .CINY1(na1678_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1680_4 ( .OUT(na1680_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na1330_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na1330_2),
                      .CINX(1'b0), .CINY1(na1678_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x17y88     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1682_2 ( .OUT(na1682_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1682_6 ( .COUTY1(na1682_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1682_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x40y86     80'h00_0078_00_0020_0C66_CA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1683_1 ( .OUT(na1683_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4407_2), .IN6(1'b1), .IN7(1'b1), .IN8(na409_1),
                      .CINX(1'b0), .CINY1(na1704_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1683_4 ( .OUT(na1683_2), .COUTY1(na1683_4), .IN1(1'b1), .IN2(na1325_1), .IN3(1'b0), .IN4(1'b0), .IN5(na4407_2), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na409_1), .CINX(1'b0), .CINY1(na1704_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x40y87     80'h00_0078_00_0020_0C66_0AC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1685_1 ( .OUT(na1685_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na410_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1683_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1685_4 ( .OUT(na1685_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na429_1), .IN5(na410_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1683_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x46y88     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1687_2 ( .OUT(na1687_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1687_6 ( .COUTY1(na1687_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1687_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x18y47     80'h00_0078_00_0020_0C66_CAC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1688_1 ( .OUT(na1688_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na173_1), .IN6(1'b1), .IN7(1'b1), .IN8(na190_2),
                      .CINX(1'b0), .CINY1(na1708_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1688_4 ( .OUT(na1688_2), .COUTY1(na1688_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na190_1), .IN5(na173_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na190_2), .CINX(1'b0), .CINY1(na1708_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x18y48     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1690_1 ( .OUT(na1690_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na192_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1688_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1690_4 ( .OUT(na1690_2), .COUTY1(na1690_4), .IN1(na192_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na192_2), .IN6(1'b1),
                      .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na1688_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x18y49     80'h00_0018_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1692_1 ( .OUT(na1692_1), .IN1(1'b1), .IN2(na193_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1690_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x30y87     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1693_2 ( .OUT(na1693_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1693_6 ( .COUTY1(na1693_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1693_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x69y85     80'h00_0078_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1694_1 ( .OUT(na1694_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na75_1), .IN7(1'b1), .IN8(na76_2),
                      .CINX(1'b0), .CINY1(na1713_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1694_4 ( .OUT(na1694_2), .COUTY1(na1694_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na76_1), .IN5(1'b1), .IN6(na75_1), .IN7(1'b1),
                      .IN8(na76_2), .CINX(1'b0), .CINY1(na1713_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x69y86     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1696_1 ( .OUT(na1696_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na78_2),
                      .CINX(1'b0), .CINY1(na1694_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1696_4 ( .OUT(na1696_2), .COUTY1(na1696_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na78_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na78_2), .CINX(1'b0), .CINY1(na1694_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x69y87     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1698_1 ( .OUT(na1698_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na79_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1696_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x64y48     80'h00_0078_00_0020_0C66_AAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1699_1 ( .OUT(na1699_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na704_2), .IN6(1'b1), .IN7(na297_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1721_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1699_4 ( .OUT(na1699_2), .COUTY1(na1699_4), .IN1(1'b1), .IN2(na2246_2), .IN3(na297_1), .IN4(1'b1), .IN5(na704_2), .IN6(1'b1),
                      .IN7(na297_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1721_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x44y83     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1701_2 ( .OUT(na1701_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1701_6 ( .COUTY1(na1701_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1701_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x47y54     80'h00_0078_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1702_1 ( .OUT(na1702_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na216_2), .IN6(1'b1), .IN7(na4302_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1727_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1702_4 ( .OUT(na1702_2), .COUTY1(na1702_4), .IN1(na216_1), .IN2(1'b1), .IN3(1'b1), .IN4(na2497_1), .IN5(na216_2), .IN6(1'b1),
                      .IN7(na4302_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na1727_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x40y85     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1704_2 ( .OUT(na1704_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1704_6 ( .COUTY1(na1704_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1704_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x30y60     80'h00_0078_00_0020_0C66_CA0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1705_1 ( .OUT(na1705_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na114_1), .IN6(1'b1), .IN7(1'b1), .IN8(na214_1),
                      .CINX(1'b0), .CINY1(na1732_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1705_4 ( .OUT(na1705_2), .COUTY1(na1705_4), .IN1(na216_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na114_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na214_1), .CINX(1'b0), .CINY1(na1732_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x30y61     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1707_1 ( .OUT(na1707_1), .IN1(na216_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1705_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x18y46     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1708_2 ( .OUT(na1708_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1708_6 ( .COUTY1(na1708_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1708_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x46y45     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1709_1 ( .OUT(na1709_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na204_2), .IN7(na201_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3234_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1709_4 ( .OUT(na1709_2), .COUTY1(na1709_4), .IN1(1'b1), .IN2(na204_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na204_2),
                      .IN7(na201_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na3234_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x46y46     80'h00_0078_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1711_1 ( .OUT(na1711_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na207_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1709_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1711_4 ( .OUT(na1711_2), .IN1(1'b1), .IN2(na207_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na207_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1709_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x69y84     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1713_2 ( .OUT(na1713_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1713_6 ( .COUTY1(na1713_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1713_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x13y50     80'h00_0078_00_0020_0C66_CC0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1714_1 ( .OUT(na1714_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na209_1), .IN7(1'b1), .IN8(na208_1),
                      .CINX(1'b0), .CINY1(na3235_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1714_4 ( .OUT(na1714_2), .COUTY1(na1714_4), .IN1(na210_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na209_1),
                      .IN7(1'b1), .IN8(na208_1), .CINX(1'b0), .CINY1(na3235_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x13y51     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1716_1 ( .OUT(na1716_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na211_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1714_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1716_4 ( .OUT(na1716_2), .IN1(1'b1), .IN2(na1353_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na211_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1714_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x56y66     80'h00_0078_00_0020_0C66_CCA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1718_1 ( .OUT(na1718_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na295_1), .IN7(1'b1), .IN8(na4171_2),
                      .CINX(1'b0), .CINY1(na3247_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1718_4 ( .OUT(na1718_2), .COUTY1(na1718_4), .IN1(1'b0), .IN2(1'b0), .IN3(na297_2), .IN4(1'b1), .IN5(1'b1), .IN6(na295_1),
                      .IN7(1'b1), .IN8(na4171_2), .CINX(1'b0), .CINY1(na3247_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x56y67     80'h00_0018_00_0010_0666_00A0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1720_1 ( .OUT(na1720_1), .IN1(1'b0), .IN2(1'b0), .IN3(na297_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1718_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x64y47     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1721_2 ( .OUT(na1721_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1721_6 ( .COUTY1(na1721_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1721_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x24y57     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1722_1 ( .OUT(na1722_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na265_2), .IN7(na264_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na3260_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1722_4 ( .OUT(na1722_2), .COUTY1(na1722_4), .IN1(1'b1), .IN2(na265_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na265_2),
                      .IN7(na264_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na3260_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x24y58     80'h00_0078_00_0020_0C66_C0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1724_1 ( .OUT(na1724_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na270_2),
                      .CINX(1'b0), .CINY1(na1722_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1724_4 ( .OUT(na1724_2), .COUTY1(na1724_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na270_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na270_2), .CINX(1'b0), .CINY1(na1722_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x24y59     80'h00_0018_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a1726_1 ( .OUT(na1726_1), .IN1(1'b1), .IN2(na268_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1724_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x47y53     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1727_2 ( .OUT(na1727_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1727_6 ( .COUTY1(na1727_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1727_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x38y62     80'h00_0078_00_0020_0C66_CAA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1728_1 ( .OUT(na1728_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1387_1), .IN6(1'b1), .IN7(1'b1), .IN8(na282_1),
                      .CINX(1'b0), .CINY1(na3267_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1728_4 ( .OUT(na1728_2), .COUTY1(na1728_4), .IN1(1'b0), .IN2(1'b0), .IN3(na283_1), .IN4(1'b1), .IN5(na1387_1), .IN6(1'b1),
                      .IN7(1'b1), .IN8(na282_1), .CINX(1'b0), .CINY1(na3267_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x38y63     80'h00_0078_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1730_1 ( .OUT(na1730_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1386_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1728_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1730_4 ( .OUT(na1730_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na284_1), .IN5(1'b1), .IN6(na1386_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1728_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x30y59     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1732_2 ( .OUT(na1732_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1732_6 ( .COUTY1(na1732_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1732_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x62y37     80'h00_0078_00_0020_0C66_CC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1733_1 ( .OUT(na1733_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na274_2), .IN7(1'b1), .IN8(na277_1),
                      .CINX(1'b0), .CINY1(na3281_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1733_4 ( .OUT(na1733_2), .COUTY1(na1733_4), .IN1(1'b1), .IN2(na274_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na274_2),
                      .IN7(1'b1), .IN8(na277_1), .CINX(1'b0), .CINY1(na3281_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x62y38     80'h00_0078_00_0020_0C66_A0A0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a1735_1 ( .OUT(na1735_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na280_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1733_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1735_4 ( .OUT(na1735_2), .IN1(1'b0), .IN2(1'b0), .IN3(na280_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na280_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1733_4), .PINX(1'b0), .PINY1(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0010_0014)) 
           _a1739 ( .GLB0(na1739_1), .GLB1(na1739_2), .GLB2(_d0), .GLB3(_d1), .CLK_FB0(_d2), .CLK_FB1(_d3), .CLK_FB2(_d4), .CLK_FB3(_d5),
                    .CLK0_0(na3222_6), .CLK0_90(na3222_5), .CLK0_180(na3222_4), .CLK0_270(na3222_3), .CLK0_BYP(1'b0), .CLK1_0(1'b0),
                    .CLK1_90(1'b0), .CLK1_180(1'b0), .CLK1_270(1'b0), .CLK1_BYP(na3229_2), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0),
                    .CLK2_270(1'b0), .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0),
                    .USR_GLB0(1'b0), .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0),
                    .USR_FB3(1'b0) );
// C_AND/D//AND/D      x53y40     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1741_1 ( .OUT(na1741_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3725_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1741_2 ( .OUT(na1741_1), .CLK(na1739_1), .EN(na1413_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1741_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1741_4 ( .OUT(na1741_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3726_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1741_5 ( .OUT(na1741_2), .CLK(na1739_1), .EN(na1413_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1741_2_i) );
// C_AND/D//AND/D      x51y38     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1743_1 ( .OUT(na1743_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3723_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1743_2 ( .OUT(na1743_1), .CLK(na1739_1), .EN(na1413_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1743_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1743_4 ( .OUT(na1743_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3724_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1743_5 ( .OUT(na1743_2), .CLK(na1739_1), .EN(na1413_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1743_2_i) );
// C_AND/D//AND/D      x57y42     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1745_1 ( .OUT(na1745_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3721_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1745_2 ( .OUT(na1745_1), .CLK(na1739_1), .EN(na1413_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1745_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1745_4 ( .OUT(na1745_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3722_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1745_5 ( .OUT(na1745_2), .CLK(na1739_1), .EN(na1413_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1745_2_i) );
// C_AND/D//AND/D      x59y42     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1747_1 ( .OUT(na1747_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3719_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1747_2 ( .OUT(na1747_1), .CLK(na1739_1), .EN(na1413_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1747_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1747_4 ( .OUT(na1747_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3720_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1747_5 ( .OUT(na1747_2), .CLK(na1739_1), .EN(na1413_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1747_2_i) );
// C_AND/D//AND/D      x35y56     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1763_1 ( .OUT(na1763_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3443_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1763_2 ( .OUT(na1763_1), .CLK(na1739_1), .EN(na1423_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1763_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1763_4 ( .OUT(na1763_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3444_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1763_5 ( .OUT(na1763_2), .CLK(na1739_1), .EN(na1423_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1763_2_i) );
// C_AND/D//AND/D      x31y56     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1765_1 ( .OUT(na1765_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3439_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1765_2 ( .OUT(na1765_1), .CLK(na1739_1), .EN(na1423_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1765_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1765_4 ( .OUT(na1765_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3442_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1765_5 ( .OUT(na1765_2), .CLK(na1739_1), .EN(na1423_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1765_2_i) );
// C_AND/D//AND/D      x45y64     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1767_1 ( .OUT(na1767_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3429_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1767_2 ( .OUT(na1767_1), .CLK(na1739_1), .EN(na1423_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1767_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1767_4 ( .OUT(na1767_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3430_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1767_5 ( .OUT(na1767_2), .CLK(na1739_1), .EN(na1423_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1767_2_i) );
// C_AND/D//AND/D      x43y60     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1769_1 ( .OUT(na1769_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3426_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1769_2 ( .OUT(na1769_1), .CLK(na1739_1), .EN(na1423_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1769_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1769_4 ( .OUT(na1769_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3427_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1769_5 ( .OUT(na1769_2), .CLK(na1739_1), .EN(na1423_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1769_2_i) );
// C_AND/D//AND/D      x41y58     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1771_1 ( .OUT(na1771_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3443_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1771_2 ( .OUT(na1771_1), .CLK(na1739_1), .EN(na1424_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1771_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1771_4 ( .OUT(na1771_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3444_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1771_5 ( .OUT(na1771_2), .CLK(na1739_1), .EN(na1424_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1771_2_i) );
// C_AND/D//AND/D      x39y58     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1773_1 ( .OUT(na1773_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3439_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1773_2 ( .OUT(na1773_1), .CLK(na1739_1), .EN(na1424_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1773_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1773_4 ( .OUT(na1773_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3442_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1773_5 ( .OUT(na1773_2), .CLK(na1739_1), .EN(na1424_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1773_2_i) );
// C_AND/D//AND/D      x39y60     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1775_1 ( .OUT(na1775_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3429_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1775_2 ( .OUT(na1775_1), .CLK(na1739_1), .EN(na1424_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1775_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1775_4 ( .OUT(na1775_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3430_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1775_5 ( .OUT(na1775_2), .CLK(na1739_1), .EN(na1424_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1775_2_i) );
// C_AND/D//AND/D      x35y54     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1777_1 ( .OUT(na1777_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3426_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1777_2 ( .OUT(na1777_1), .CLK(na1739_1), .EN(na1424_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1777_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1777_4 ( .OUT(na1777_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3427_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1777_5 ( .OUT(na1777_2), .CLK(na1739_1), .EN(na1424_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1777_2_i) );
// C_AND/D//AND/D      x48y68     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1780_1 ( .OUT(na1780_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3423_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1780_2 ( .OUT(na1780_1), .CLK(na1739_1), .EN(na1420_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1780_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1780_4 ( .OUT(na1780_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3424_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1780_5 ( .OUT(na1780_2), .CLK(na1739_1), .EN(na1420_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1780_2_i) );
// C_AND/D//AND/D      x44y66     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1782_1 ( .OUT(na1782_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3420_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1782_2 ( .OUT(na1782_1), .CLK(na1739_1), .EN(na1420_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1782_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1782_4 ( .OUT(na1782_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3421_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1782_5 ( .OUT(na1782_2), .CLK(na1739_1), .EN(na1420_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1782_2_i) );
// C_AND/D//AND/D      x46y74     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1784_1 ( .OUT(na1784_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3416_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1784_2 ( .OUT(na1784_1), .CLK(na1739_1), .EN(na1420_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1784_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1784_4 ( .OUT(na1784_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3417_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1784_5 ( .OUT(na1784_2), .CLK(na1739_1), .EN(na1420_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1784_2_i) );
// C_AND/D//AND/D      x46y76     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1786_1 ( .OUT(na1786_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3413_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1786_2 ( .OUT(na1786_1), .CLK(na1739_1), .EN(na1420_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1786_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1786_4 ( .OUT(na1786_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3414_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1786_5 ( .OUT(na1786_2), .CLK(na1739_1), .EN(na1420_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1786_2_i) );
// C_AND/D//AND/D      x48y66     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1788_1 ( .OUT(na1788_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3423_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1788_2 ( .OUT(na1788_1), .CLK(na1739_1), .EN(na1421_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1788_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1788_4 ( .OUT(na1788_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3424_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1788_5 ( .OUT(na1788_2), .CLK(na1739_1), .EN(na1421_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1788_2_i) );
// C_AND/D//AND/D      x46y70     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1790_1 ( .OUT(na1790_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3420_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1790_2 ( .OUT(na1790_1), .CLK(na1739_1), .EN(na1421_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1790_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1790_4 ( .OUT(na1790_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3421_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1790_5 ( .OUT(na1790_2), .CLK(na1739_1), .EN(na1421_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1790_2_i) );
// C_AND/D//AND/D      x48y72     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1792_1 ( .OUT(na1792_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3416_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1792_2 ( .OUT(na1792_1), .CLK(na1739_1), .EN(na1421_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1792_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1792_4 ( .OUT(na1792_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3417_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1792_5 ( .OUT(na1792_2), .CLK(na1739_1), .EN(na1421_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1792_2_i) );
// C_AND/D//AND/D      x46y66     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1794_1 ( .OUT(na1794_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3413_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1794_2 ( .OUT(na1794_1), .CLK(na1739_1), .EN(na1421_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1794_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1794_4 ( .OUT(na1794_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3414_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1794_5 ( .OUT(na1794_2), .CLK(na1739_1), .EN(na1421_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1794_2_i) );
// C_AND/D//AND/D      x40y43     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1811_1 ( .OUT(na1811_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3531_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1811_2 ( .OUT(na1811_1), .CLK(na1739_1), .EN(na1417_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1811_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1811_4 ( .OUT(na1811_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3532_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1811_5 ( .OUT(na1811_2), .CLK(na1739_1), .EN(na1417_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1811_2_i) );
// C_AND/D//AND/D      x38y43     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1813_1 ( .OUT(na1813_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3529_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1813_2 ( .OUT(na1813_1), .CLK(na1739_1), .EN(na1417_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1813_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1813_4 ( .OUT(na1813_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1813_5 ( .OUT(na1813_2), .CLK(na1739_1), .EN(na1417_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1813_2_i) );
// C_AND/D//AND/D      x36y45     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1815_1 ( .OUT(na1815_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3527_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1815_2 ( .OUT(na1815_1), .CLK(na1739_1), .EN(na1417_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1815_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1815_4 ( .OUT(na1815_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3528_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1815_5 ( .OUT(na1815_2), .CLK(na1739_1), .EN(na1417_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1815_2_i) );
// C_AND/D//AND/D      x38y39     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1817_1 ( .OUT(na1817_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3525_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1817_2 ( .OUT(na1817_1), .CLK(na1739_1), .EN(na1417_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1817_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1817_4 ( .OUT(na1817_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3526_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1817_5 ( .OUT(na1817_2), .CLK(na1739_1), .EN(na1417_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1817_2_i) );
// C_AND/D//AND/D      x26y39     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1819_1 ( .OUT(na1819_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3531_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1819_2 ( .OUT(na1819_1), .CLK(na1739_1), .EN(na1416_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1819_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1819_4 ( .OUT(na1819_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3532_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1819_5 ( .OUT(na1819_2), .CLK(na1739_1), .EN(na1416_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1819_2_i) );
// C_AND/D//AND/D      x24y39     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1821_1 ( .OUT(na1821_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3529_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1821_2 ( .OUT(na1821_1), .CLK(na1739_1), .EN(na1416_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1821_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1821_4 ( .OUT(na1821_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1821_5 ( .OUT(na1821_2), .CLK(na1739_1), .EN(na1416_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1821_2_i) );
// C_AND/D//AND/D      x40y45     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1823_1 ( .OUT(na1823_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3527_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1823_2 ( .OUT(na1823_1), .CLK(na1739_1), .EN(na1416_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1823_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1823_4 ( .OUT(na1823_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3528_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1823_5 ( .OUT(na1823_2), .CLK(na1739_1), .EN(na1416_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1823_2_i) );
// C_AND/D//AND/D      x38y47     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1825_1 ( .OUT(na1825_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3525_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1825_2 ( .OUT(na1825_1), .CLK(na1739_1), .EN(na1416_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1825_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1825_4 ( .OUT(na1825_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3526_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1825_5 ( .OUT(na1825_2), .CLK(na1739_1), .EN(na1416_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1825_2_i) );
// C_AND/D//AND/D      x56y49     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1862_1 ( .OUT(na1862_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3717_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1862_2 ( .OUT(na1862_1), .CLK(na1739_1), .EN(na1411_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1862_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1862_4 ( .OUT(na1862_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3718_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1862_5 ( .OUT(na1862_2), .CLK(na1739_1), .EN(na1411_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1862_2_i) );
// C_AND/D//AND/D      x58y49     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1864_1 ( .OUT(na1864_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3715_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1864_2 ( .OUT(na1864_1), .CLK(na1739_1), .EN(na1411_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1864_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1864_4 ( .OUT(na1864_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3716_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1864_5 ( .OUT(na1864_2), .CLK(na1739_1), .EN(na1411_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1864_2_i) );
// C_AND/D//AND/D      x58y53     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1866_1 ( .OUT(na1866_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3713_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1866_2 ( .OUT(na1866_1), .CLK(na1739_1), .EN(na1411_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1866_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1866_4 ( .OUT(na1866_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3714_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1866_5 ( .OUT(na1866_2), .CLK(na1739_1), .EN(na1411_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1866_2_i) );
// C_AND/D//AND/D      x54y47     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1868_1 ( .OUT(na1868_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3711_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1868_2 ( .OUT(na1868_1), .CLK(na1739_1), .EN(na1411_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1868_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1868_4 ( .OUT(na1868_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3712_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1868_5 ( .OUT(na1868_2), .CLK(na1739_1), .EN(na1411_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1868_2_i) );
// C_AND/D//AND/D      x59y40     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1878_1 ( .OUT(na1878_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3725_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1878_2 ( .OUT(na1878_1), .CLK(na1739_1), .EN(na1414_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1878_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1878_4 ( .OUT(na1878_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3726_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1878_5 ( .OUT(na1878_2), .CLK(na1739_1), .EN(na1414_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1878_2_i) );
// C_AND/D//AND/D      x57y38     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1880_1 ( .OUT(na1880_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3723_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1880_2 ( .OUT(na1880_1), .CLK(na1739_1), .EN(na1414_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1880_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1880_4 ( .OUT(na1880_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3724_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1880_5 ( .OUT(na1880_2), .CLK(na1739_1), .EN(na1414_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1880_2_i) );
// C_AND/D//AND/D      x57y40     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1882_1 ( .OUT(na1882_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3721_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1882_2 ( .OUT(na1882_1), .CLK(na1739_1), .EN(na1414_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1882_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1882_4 ( .OUT(na1882_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3722_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1882_5 ( .OUT(na1882_2), .CLK(na1739_1), .EN(na1414_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1882_2_i) );
// C_AND/D//AND/D      x55y40     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1884_1 ( .OUT(na1884_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3719_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1884_2 ( .OUT(na1884_1), .CLK(na1739_1), .EN(na1414_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1884_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1884_4 ( .OUT(na1884_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3720_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1884_5 ( .OUT(na1884_2), .CLK(na1739_1), .EN(na1414_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1884_2_i) );
// C_AND/D//AND/D      x51y49     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1887_1 ( .OUT(na1887_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3717_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1887_2 ( .OUT(na1887_1), .CLK(na1739_1), .EN(na1410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1887_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1887_4 ( .OUT(na1887_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3718_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1887_5 ( .OUT(na1887_2), .CLK(na1739_1), .EN(na1410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1887_2_i) );
// C_AND/D//AND/D      x52y47     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1889_1 ( .OUT(na1889_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3715_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1889_2 ( .OUT(na1889_1), .CLK(na1739_1), .EN(na1410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1889_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1889_4 ( .OUT(na1889_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3716_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1889_5 ( .OUT(na1889_2), .CLK(na1739_1), .EN(na1410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1889_2_i) );
// C_AND/D//AND/D      x60y55     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1891_1 ( .OUT(na1891_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3713_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1891_2 ( .OUT(na1891_1), .CLK(na1739_1), .EN(na1410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1891_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1891_4 ( .OUT(na1891_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3714_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1891_5 ( .OUT(na1891_2), .CLK(na1739_1), .EN(na1410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1891_2_i) );
// C_AND/D//AND/D      x60y53     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1893_1 ( .OUT(na1893_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3711_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1893_2 ( .OUT(na1893_1), .CLK(na1739_1), .EN(na1410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1893_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1893_4 ( .OUT(na1893_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3712_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1893_5 ( .OUT(na1893_2), .CLK(na1739_1), .EN(na1410_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na1893_2_i) );
// C_///AND/D      x52y60     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1984_4 ( .OUT(na1984_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3712_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1984_5 ( .OUT(na1984_2), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1984_2_i) );
// C_AND/D///      x66y66     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1985_1 ( .OUT(na1985_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1891_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1985_2 ( .OUT(na1985_1), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1985_1_i) );
// C_AND/D//AND/D      x65y68     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1986_1 ( .OUT(na1986_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1891_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1986_2 ( .OUT(na1986_1), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1986_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1986_4 ( .OUT(na1986_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1893_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1986_5 ( .OUT(na1986_2), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1986_2_i) );
// C_///AND/D      x61y66     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1989_4 ( .OUT(na1989_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2120_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1989_5 ( .OUT(na1989_2), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1989_2_i) );
// C_AND/D//AND/D      x62y70     80'h00_FA00_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1990_1 ( .OUT(na1990_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2122_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1990_2 ( .OUT(na1990_1), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1990_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1990_4 ( .OUT(na1990_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2120_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1990_5 ( .OUT(na1990_2), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1990_2_i) );
// C_AND/D///      x62y65     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1991_1 ( .OUT(na1991_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2122_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1991_2 ( .OUT(na1991_1), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1991_1_i) );
// C_AND/D//AND/D      x61y68     80'h00_FA00_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1993_1 ( .OUT(na1993_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3711_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1993_2 ( .OUT(na1993_1), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1993_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1993_4 ( .OUT(na1993_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2124_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1993_5 ( .OUT(na1993_2), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1993_2_i) );
// C_///AND/D      x59y54     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1994_4 ( .OUT(na1994_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1866_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1994_5 ( .OUT(na1994_2), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1994_2_i) );
// C_AND/D///      x55y54     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1995_1 ( .OUT(na1995_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1866_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1995_2 ( .OUT(na1995_1), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1995_1_i) );
// C_///AND/D      x53y52     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1996_4 ( .OUT(na1996_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1868_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1996_5 ( .OUT(na1996_2), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1996_2_i) );
// C_AND/D///      x53y52     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1997_1 ( .OUT(na1997_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1868_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1997_2 ( .OUT(na1997_1), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1997_1_i) );
// C_///AND/D      x43y48     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1998_4 ( .OUT(na1998_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3718_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1998_5 ( .OUT(na1998_2), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1998_2_i) );
// C_AND/D///      x54y57     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1999_1 ( .OUT(na1999_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2124_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1999_2 ( .OUT(na1999_1), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1999_1_i) );
// C_///AND/D      x50y52     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2000_4 ( .OUT(na2000_2_i), .IN1(na1887_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2000_5 ( .OUT(na2000_2), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2000_2_i) );
// C_AND/D//AND/D      x49y51     80'h00_FA00_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2001_1 ( .OUT(na2001_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1887_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2001_2 ( .OUT(na2001_1), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2001_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2001_4 ( .OUT(na2001_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1889_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2001_5 ( .OUT(na2001_2), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2001_2_i) );
// C_AND/D///      x50y51     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2002_1 ( .OUT(na2002_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1889_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2002_2 ( .OUT(na2002_1), .CLK(na1739_1), .EN(na54_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2002_1_i) );
// C_AND/D//AND/D      x66y76     80'h00_F600_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2011_1 ( .OUT(na2011_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2011_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2011_2 ( .OUT(na2011_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2011_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2011_4 ( .OUT(na2011_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2013_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2011_5 ( .OUT(na2011_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2011_2_i) );
// C_AND/D//AND/D      x60y65     80'h00_F600_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2013_1 ( .OUT(na2013_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2013_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2013_2 ( .OUT(na2013_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2013_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2013_4 ( .OUT(na2013_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2015_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2013_5 ( .OUT(na2013_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2013_2_i) );
// C_AND/D//AND/D      x50y60     80'h00_F600_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2015_1 ( .OUT(na2015_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2015_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2015_2 ( .OUT(na2015_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2015_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2015_4 ( .OUT(na2015_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2017_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2015_5 ( .OUT(na2015_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2015_2_i) );
// C_AND/D//AND/D      x44y55     80'h00_F600_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2017_1 ( .OUT(na2017_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2017_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2017_2 ( .OUT(na2017_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2017_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2017_4 ( .OUT(na2017_2_i), .IN1(na2019_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2017_5 ( .OUT(na2017_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2017_2_i) );
// C_AND/D//AND/D      x21y57     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2019_1 ( .OUT(na2019_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2019_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2019_2 ( .OUT(na2019_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2019_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2019_4 ( .OUT(na2019_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2021_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2019_5 ( .OUT(na2019_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2019_2_i) );
// C_AND/D//AND/D      x16y47     80'h00_F600_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2021_1 ( .OUT(na2021_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2021_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2021_2 ( .OUT(na2021_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2021_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2021_4 ( .OUT(na2021_2_i), .IN1(na2023_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2021_5 ( .OUT(na2021_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2021_2_i) );
// C_AND/D//AND/D      x13y45     80'h00_F600_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2023_1 ( .OUT(na2023_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2023_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2023_2 ( .OUT(na2023_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2023_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2023_4 ( .OUT(na2023_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2025_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2023_5 ( .OUT(na2023_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2023_2_i) );
// C_AND/D//AND/D      x14y44     80'h00_F600_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2025_1 ( .OUT(na2025_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2025_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2025_2 ( .OUT(na2025_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2025_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2025_4 ( .OUT(na2025_2_i), .IN1(1'b1), .IN2(na2027_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2025_5 ( .OUT(na2025_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2025_2_i) );
// C_AND/D//AND/D      x15y40     80'h00_F600_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2027_1 ( .OUT(na2027_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2027_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2027_2 ( .OUT(na2027_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2027_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2027_4 ( .OUT(na2027_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2029_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2027_5 ( .OUT(na2027_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2027_2_i) );
// C_AND/D//AND/D      x14y39     80'h00_F600_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2029_1 ( .OUT(na2029_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2029_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2029_2 ( .OUT(na2029_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2029_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2029_4 ( .OUT(na2029_2_i), .IN1(na2031_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2029_5 ( .OUT(na2029_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2029_2_i) );
// C_AND/D//AND/D      x13y37     80'h00_F600_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2031_1 ( .OUT(na2031_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2031_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2031_2 ( .OUT(na2031_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2031_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2031_4 ( .OUT(na2031_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2033_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2031_5 ( .OUT(na2031_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2031_2_i) );
// C_AND/D//AND/D      x14y42     80'h00_F600_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2033_1 ( .OUT(na2033_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2033_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2033_2 ( .OUT(na2033_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2033_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2033_4 ( .OUT(na2033_2_i), .IN1(na2035_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2033_5 ( .OUT(na2033_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2033_2_i) );
// C_AND/D//AND/D      x15y45     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2035_1 ( .OUT(na2035_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2035_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2035_2 ( .OUT(na2035_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2035_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2035_4 ( .OUT(na2035_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2037_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2035_5 ( .OUT(na2035_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2035_2_i) );
// C_AND/D//AND/D      x24y61     80'h00_F600_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2037_1 ( .OUT(na2037_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2037_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2037_2 ( .OUT(na2037_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2037_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2037_4 ( .OUT(na2037_2_i), .IN1(na2039_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2037_5 ( .OUT(na2037_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2037_2_i) );
// C_AND/D//AND/D      x47y57     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2039_1 ( .OUT(na2039_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2039_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2039_2 ( .OUT(na2039_1), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2039_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2039_4 ( .OUT(na2039_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2041_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2039_5 ( .OUT(na2039_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2039_2_i) );
// C_///AND/D      x62y61     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2041_4 ( .OUT(na2041_2_i), .IN1(na525_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2041_5 ( .OUT(na2041_2), .CLK(na1739_1), .EN(~na1431_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2041_2_i) );
// C_AND/D//AND/D      x69y83     80'h00_FA00_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2091_1 ( .OUT(na2091_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2091_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2091_2 ( .OUT(na2091_1), .CLK(na1739_1), .EN(na1435_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2091_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2091_4 ( .OUT(na2091_2_i), .IN1(1'b1), .IN2(na2093_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2091_5 ( .OUT(na2091_2), .CLK(na1739_1), .EN(na1435_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2091_2_i) );
// C_AND/D///      x69y82     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2093_1 ( .OUT(na2093_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na534_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2093_2 ( .OUT(na2093_1), .CLK(na1739_1), .EN(na1435_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2093_1_i) );
// C_AND/D//AND/D      x50y41     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2118_1 ( .OUT(na2118_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3717_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2118_2 ( .OUT(na2118_1), .CLK(na1739_1), .EN(na1409_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2118_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2118_4 ( .OUT(na2118_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3718_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2118_5 ( .OUT(na2118_2), .CLK(na1739_1), .EN(na1409_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2118_2_i) );
// C_AND/D//AND/D      x52y51     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2120_1 ( .OUT(na2120_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3715_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2120_2 ( .OUT(na2120_1), .CLK(na1739_1), .EN(na1409_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2120_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2120_4 ( .OUT(na2120_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3716_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2120_5 ( .OUT(na2120_2), .CLK(na1739_1), .EN(na1409_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2120_2_i) );
// C_AND/D//AND/D      x51y51     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2122_1 ( .OUT(na2122_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3713_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2122_2 ( .OUT(na2122_1), .CLK(na1739_1), .EN(na1409_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2122_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2122_4 ( .OUT(na2122_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3714_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2122_5 ( .OUT(na2122_2), .CLK(na1739_1), .EN(na1409_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2122_2_i) );
// C_AND/D//AND/D      x54y55     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2124_1 ( .OUT(na2124_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3711_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2124_2 ( .OUT(na2124_1), .CLK(na1739_1), .EN(na1409_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2124_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2124_4 ( .OUT(na2124_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3712_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2124_5 ( .OUT(na2124_2), .CLK(na1739_1), .EN(na1409_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2124_2_i) );
// C_AND/D//AND/D      x69y58     80'h00_FE00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2125_1 ( .OUT(na2125_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2125_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2125_2 ( .OUT(na2125_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2125_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2125_4 ( .OUT(na2125_2_i), .IN1(1'b1), .IN2(na2127_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2125_5 ( .OUT(na2125_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2125_2_i) );
// C_AND/D//AND/D      x69y60     80'h00_FE00_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2127_1 ( .OUT(na2127_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2127_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2127_2 ( .OUT(na2127_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2127_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2127_4 ( .OUT(na2127_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2129_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2127_5 ( .OUT(na2127_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2127_2_i) );
// C_AND/D//AND/D      x70y63     80'h00_FE00_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2129_1 ( .OUT(na2129_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2129_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2129_2 ( .OUT(na2129_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2129_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2129_4 ( .OUT(na2129_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na597_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2129_5 ( .OUT(na2129_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2129_2_i) );
// C_///AND/D      x58y40     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2221_4 ( .OUT(na2221_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3720_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2221_5 ( .OUT(na2221_2), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2221_2_i) );
// C_AND/D///      x67y53     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2222_1 ( .OUT(na2222_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1745_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2222_2 ( .OUT(na2222_1), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2222_1_i) );
// C_AND/D//AND/D      x68y51     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2223_1 ( .OUT(na2223_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1745_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2223_2 ( .OUT(na2223_1), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2223_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2223_4 ( .OUT(na2223_2_i), .IN1(1'b1), .IN2(na1747_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2223_5 ( .OUT(na2223_2), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2223_2_i) );
// C_///AND/D      x60y61     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2226_4 ( .OUT(na2226_2_i), .IN1(1'b1), .IN2(na2354_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2226_5 ( .OUT(na2226_2), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2226_2_i) );
// C_AND/D//AND/D      x55y60     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2228_1 ( .OUT(na2228_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2356_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2228_2 ( .OUT(na2228_1), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2228_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2228_4 ( .OUT(na2228_2_i), .IN1(1'b1), .IN2(na2356_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2228_5 ( .OUT(na2228_2), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2228_2_i) );
// C_AND/D//AND/D      x57y59     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2229_1 ( .OUT(na2229_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2358_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2229_2 ( .OUT(na2229_1), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2229_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2229_4 ( .OUT(na2229_2_i), .IN1(1'b1), .IN2(na2354_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2229_5 ( .OUT(na2229_2), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2229_2_i) );
// C_AND/D///      x52y50     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2230_1 ( .OUT(na2230_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3719_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2230_2 ( .OUT(na2230_1), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2230_1_i) );
// C_AND/D///      x61y42     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2231_1 ( .OUT(na2231_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1882_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2231_2 ( .OUT(na2231_1), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2231_1_i) );
// C_AND/D///      x55y42     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2232_1 ( .OUT(na2232_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1882_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2232_2 ( .OUT(na2232_1), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2232_1_i) );
// C_///AND/D      x61y40     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2233_4 ( .OUT(na2233_2_i), .IN1(1'b1), .IN2(na1884_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2233_5 ( .OUT(na2233_2), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2233_2_i) );
// C_AND/D///      x55y38     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2234_1 ( .OUT(na2234_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1884_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2234_2 ( .OUT(na2234_1), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2234_1_i) );
// C_///AND/D      x43y40     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2235_4 ( .OUT(na2235_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3726_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2235_5 ( .OUT(na2235_2), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2235_2_i) );
// C_AND/D///      x52y44     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2236_1 ( .OUT(na2236_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2358_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2236_2 ( .OUT(na2236_1), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2236_1_i) );
// C_///AND/D      x56y40     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2237_4 ( .OUT(na2237_2_i), .IN1(1'b1), .IN2(na1741_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2237_5 ( .OUT(na2237_2), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2237_2_i) );
// C_AND/D//AND/D      x53y44     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2238_1 ( .OUT(na2238_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1741_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2238_2 ( .OUT(na2238_1), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2238_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2238_4 ( .OUT(na2238_2_i), .IN1(1'b1), .IN2(na1743_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2238_5 ( .OUT(na2238_2), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2238_2_i) );
// C_AND/D///      x52y41     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2239_1 ( .OUT(na2239_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1743_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2239_2 ( .OUT(na2239_1), .CLK(na1739_1), .EN(na275_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2239_1_i) );
// C_///AND/D      x65y48     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2246_4 ( .OUT(na2246_2_i), .IN1(na704_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2246_5 ( .OUT(na2246_2), .CLK(na1739_1), .EN(na1458_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2246_2_i) );
// C_AND/D//AND/D      x57y62     80'h00_F600_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2248_1 ( .OUT(na2248_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2248_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2248_2 ( .OUT(na2248_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2248_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2248_4 ( .OUT(na2248_2_i), .IN1(na2250_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2248_5 ( .OUT(na2248_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2248_2_i) );
// C_AND/D//AND/D      x49y55     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2250_1 ( .OUT(na2250_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2250_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2250_2 ( .OUT(na2250_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2250_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2250_4 ( .OUT(na2250_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2252_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2250_5 ( .OUT(na2250_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2250_2_i) );
// C_AND/D//AND/D      x46y53     80'h00_F600_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2252_1 ( .OUT(na2252_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2252_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2252_2 ( .OUT(na2252_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2252_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2252_4 ( .OUT(na2252_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2254_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2252_5 ( .OUT(na2252_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2252_2_i) );
// C_AND/D//AND/D      x38y52     80'h00_F600_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2254_1 ( .OUT(na2254_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2254_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2254_2 ( .OUT(na2254_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2254_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2254_4 ( .OUT(na2254_2_i), .IN1(na2256_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2254_5 ( .OUT(na2254_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2254_2_i) );
// C_AND/D//AND/D      x19y41     80'h00_F600_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2256_1 ( .OUT(na2256_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2256_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2256_2 ( .OUT(na2256_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2256_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2256_4 ( .OUT(na2256_2_i), .IN1(na2258_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2256_5 ( .OUT(na2256_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2256_2_i) );
// C_AND/D//AND/D      x19y39     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2258_1 ( .OUT(na2258_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2258_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2258_2 ( .OUT(na2258_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2258_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2258_4 ( .OUT(na2258_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2260_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2258_5 ( .OUT(na2258_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2258_2_i) );
// C_AND/D//AND/D      x16y39     80'h00_F600_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2260_1 ( .OUT(na2260_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2260_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2260_2 ( .OUT(na2260_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2260_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2260_4 ( .OUT(na2260_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2262_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2260_5 ( .OUT(na2260_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2260_2_i) );
// C_AND/D//AND/D      x16y38     80'h00_F600_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2262_1 ( .OUT(na2262_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2262_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2262_2 ( .OUT(na2262_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2262_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2262_4 ( .OUT(na2262_2_i), .IN1(na2264_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2262_5 ( .OUT(na2262_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2262_2_i) );
// C_AND/D//AND/D      x15y37     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2264_1 ( .OUT(na2264_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2264_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2264_2 ( .OUT(na2264_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2264_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2264_4 ( .OUT(na2264_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2266_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2264_5 ( .OUT(na2264_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2264_2_i) );
// C_AND/D//AND/D      x16y35     80'h00_F600_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2266_1 ( .OUT(na2266_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2266_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2266_2 ( .OUT(na2266_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2266_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2266_4 ( .OUT(na2266_2_i), .IN1(1'b1), .IN2(na2268_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2266_5 ( .OUT(na2266_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2266_2_i) );
// C_AND/D//AND/D      x15y38     80'h00_F600_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2268_1 ( .OUT(na2268_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2268_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2268_2 ( .OUT(na2268_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2268_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2268_4 ( .OUT(na2268_2_i), .IN1(na2270_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2268_5 ( .OUT(na2268_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2268_2_i) );
// C_AND/D//AND/D      x15y39     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2270_1 ( .OUT(na2270_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2270_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2270_2 ( .OUT(na2270_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2270_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2270_4 ( .OUT(na2270_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2272_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2270_5 ( .OUT(na2270_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2270_2_i) );
// C_AND/D//AND/D      x16y43     80'h00_F600_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2272_1 ( .OUT(na2272_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2272_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2272_2 ( .OUT(na2272_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2272_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2272_4 ( .OUT(na2272_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2274_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2272_5 ( .OUT(na2272_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2272_2_i) );
// C_AND/D//AND/D      x16y46     80'h00_F600_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2274_1 ( .OUT(na2274_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2274_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2274_2 ( .OUT(na2274_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2274_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2274_4 ( .OUT(na2274_2_i), .IN1(na2276_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2274_5 ( .OUT(na2274_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2274_2_i) );
// C_AND/D//AND/D      x31y49     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2276_1 ( .OUT(na2276_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2276_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2276_2 ( .OUT(na2276_1), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2276_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2276_4 ( .OUT(na2276_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2278_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2276_5 ( .OUT(na2276_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2276_2_i) );
// C_///AND/D      x48y51     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2278_4 ( .OUT(na2278_2_i), .IN1(na709_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2278_5 ( .OUT(na2278_2), .CLK(na1739_1), .EN(~na1453_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2278_2_i) );
// C_AND/D//AND/D      x32y62     80'h00_FA00_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2337_1 ( .OUT(na2337_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2337_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2337_2 ( .OUT(na2337_1), .CLK(na1739_1), .EN(na1457_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2337_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2337_4 ( .OUT(na2337_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2339_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2337_5 ( .OUT(na2337_2), .CLK(na1739_1), .EN(na1457_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2337_2_i) );
// C_AND/D///      x42y57     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2339_1 ( .OUT(na2339_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na713_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2339_2 ( .OUT(na2339_1), .CLK(na1739_1), .EN(na1457_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2339_1_i) );
// C_///AND/D      x67y66     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2350_4 ( .OUT(na2350_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na519_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2350_5 ( .OUT(na2350_2), .CLK(na1739_1), .EN(na1437_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2350_2_i) );
// C_AND/D//AND/D      x49y38     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2352_1 ( .OUT(na2352_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3725_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2352_2 ( .OUT(na2352_1), .CLK(na1739_1), .EN(na1412_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2352_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2352_4 ( .OUT(na2352_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3726_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2352_5 ( .OUT(na2352_2), .CLK(na1739_1), .EN(na1412_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2352_2_i) );
// C_AND/D//AND/D      x53y42     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2354_1 ( .OUT(na2354_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3723_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2354_2 ( .OUT(na2354_1), .CLK(na1739_1), .EN(na1412_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2354_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2354_4 ( .OUT(na2354_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3724_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2354_5 ( .OUT(na2354_2), .CLK(na1739_1), .EN(na1412_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2354_2_i) );
// C_AND/D//AND/D      x51y42     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2356_1 ( .OUT(na2356_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3721_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2356_2 ( .OUT(na2356_1), .CLK(na1739_1), .EN(na1412_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2356_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2356_4 ( .OUT(na2356_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3722_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2356_5 ( .OUT(na2356_2), .CLK(na1739_1), .EN(na1412_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2356_2_i) );
// C_AND/D//AND/D      x53y46     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2358_1 ( .OUT(na2358_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3719_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2358_2 ( .OUT(na2358_1), .CLK(na1739_1), .EN(na1412_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2358_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2358_4 ( .OUT(na2358_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3720_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2358_5 ( .OUT(na2358_2), .CLK(na1739_1), .EN(na1412_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2358_2_i) );
// C_AND/D//AND/D      x69y42     80'h00_FE00_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2359_1 ( .OUT(na2359_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2359_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2359_2 ( .OUT(na2359_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2359_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2359_4 ( .OUT(na2359_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2361_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2359_5 ( .OUT(na2359_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2359_2_i) );
// C_AND/D//AND/D      x68y41     80'h00_FE00_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2361_1 ( .OUT(na2361_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2361_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2361_2 ( .OUT(na2361_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2361_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2361_4 ( .OUT(na2361_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2363_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2361_5 ( .OUT(na2361_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2361_2_i) );
// C_AND/D//AND/D      x66y44     80'h00_FE00_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2363_1 ( .OUT(na2363_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2363_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2363_2 ( .OUT(na2363_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2363_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2363_4 ( .OUT(na2363_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na784_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2363_5 ( .OUT(na2363_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2363_2_i) );
// C_AND/D///      x25y41     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2472_1 ( .OUT(na2472_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3526_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2472_2 ( .OUT(na2472_1), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2472_1_i) );
// C_///AND/D      x34y60     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2473_4 ( .OUT(na2473_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1823_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2473_5 ( .OUT(na2473_2), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2473_2_i) );
// C_AND/D//AND/D      x29y58     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2474_1 ( .OUT(na2474_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1823_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2474_2 ( .OUT(na2474_1), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2474_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2474_4 ( .OUT(na2474_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1825_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2474_5 ( .OUT(na2474_2), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2474_2_i) );
// C_AND/D///      x19y52     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2477_1 ( .OUT(na2477_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2595_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2477_2 ( .OUT(na2477_1), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2477_1_i) );
// C_AND/D//AND/D      x19y56     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2478_1 ( .OUT(na2478_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2597_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2478_2 ( .OUT(na2478_1), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2478_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2478_4 ( .OUT(na2478_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2595_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2478_5 ( .OUT(na2478_2), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2478_2_i) );
// C_///AND/D      x19y51     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2479_4 ( .OUT(na2479_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2597_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2479_5 ( .OUT(na2479_2), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2479_2_i) );
// C_AND/D//AND/D      x20y49     80'h00_FA00_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2481_1 ( .OUT(na2481_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3525_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2481_2 ( .OUT(na2481_1), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2481_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2481_4 ( .OUT(na2481_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2599_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2481_5 ( .OUT(na2481_2), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2481_2_i) );
// C_AND/D///      x29y44     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2482_1 ( .OUT(na2482_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1815_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2482_2 ( .OUT(na2482_1), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2482_1_i) );
// C_///AND/D      x26y46     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2483_4 ( .OUT(na2483_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1815_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2483_5 ( .OUT(na2483_2), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2483_2_i) );
// C_AND/D///      x38y45     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2484_1 ( .OUT(na2484_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1817_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2484_2 ( .OUT(na2484_1), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2484_1_i) );
// C_///AND/D      x35y38     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2485_4 ( .OUT(na2485_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1817_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2485_5 ( .OUT(na2485_2), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2485_2_i) );
// C_AND/D///      x35y38     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2486_1 ( .OUT(na2486_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3532_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2486_2 ( .OUT(na2486_1), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2486_1_i) );
// C_///AND/D      x20y45     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2487_4 ( .OUT(na2487_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2599_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2487_5 ( .OUT(na2487_2), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2487_2_i) );
// C_AND/D///      x22y43     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2488_1 ( .OUT(na2488_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1819_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2488_2 ( .OUT(na2488_1), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2488_1_i) );
// C_AND/D//AND/D      x22y44     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2489_1 ( .OUT(na2489_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1819_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2489_2 ( .OUT(na2489_1), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2489_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2489_4 ( .OUT(na2489_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1821_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2489_5 ( .OUT(na2489_2), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2489_2_i) );
// C_///AND/D      x13y39     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2490_4 ( .OUT(na2490_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1821_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2490_5 ( .OUT(na2490_2), .CLK(na1739_1), .EN(na121_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2490_2_i) );
// C_AND/D///      x38y50     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2497_1 ( .OUT(na2497_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na881_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2497_2 ( .OUT(na2497_1), .CLK(na1739_1), .EN(na1480_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2497_1_i) );
// C_AND/D//AND/D      x18y52     80'h00_F600_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2499_1 ( .OUT(na2499_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2499_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2499_2 ( .OUT(na2499_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2499_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2499_4 ( .OUT(na2499_2_i), .IN1(na2501_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2499_5 ( .OUT(na2499_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2499_2_i) );
// C_AND/D//AND/D      x15y43     80'h00_F600_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2501_1 ( .OUT(na2501_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2501_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2501_2 ( .OUT(na2501_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2501_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2501_4 ( .OUT(na2501_2_i), .IN1(1'b1), .IN2(na2503_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2501_5 ( .OUT(na2501_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2501_2_i) );
// C_AND/D//AND/D      x15y44     80'h00_F600_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2503_1 ( .OUT(na2503_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2503_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2503_2 ( .OUT(na2503_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2503_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2503_4 ( .OUT(na2503_2_i), .IN1(na2505_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2503_5 ( .OUT(na2503_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2503_2_i) );
// C_AND/D//AND/D      x13y41     80'h00_F600_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2505_1 ( .OUT(na2505_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2505_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2505_2 ( .OUT(na2505_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2505_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2505_4 ( .OUT(na2505_2_i), .IN1(1'b1), .IN2(na2507_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2505_5 ( .OUT(na2505_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2505_2_i) );
// C_AND/D//AND/D      x15y42     80'h00_F600_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2507_1 ( .OUT(na2507_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2507_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2507_2 ( .OUT(na2507_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2507_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2507_4 ( .OUT(na2507_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2509_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2507_5 ( .OUT(na2507_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2507_2_i) );
// C_AND/D//AND/D      x18y39     80'h00_F600_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2509_1 ( .OUT(na2509_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2509_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2509_2 ( .OUT(na2509_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2509_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2509_4 ( .OUT(na2509_2_i), .IN1(1'b1), .IN2(na2511_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2509_5 ( .OUT(na2509_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2509_2_i) );
// C_AND/D//AND/D      x17y38     80'h00_F600_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2511_1 ( .OUT(na2511_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2511_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2511_2 ( .OUT(na2511_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2511_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2511_4 ( .OUT(na2511_2_i), .IN1(na2513_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2511_5 ( .OUT(na2511_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2511_2_i) );
// C_AND/D//AND/D      x17y37     80'h00_F600_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2513_1 ( .OUT(na2513_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2513_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2513_2 ( .OUT(na2513_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2513_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2513_4 ( .OUT(na2513_2_i), .IN1(1'b1), .IN2(na2515_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2513_5 ( .OUT(na2513_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2513_2_i) );
// C_AND/D//AND/D      x19y38     80'h00_F600_80_0000_0C88_FCCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2515_1 ( .OUT(na2515_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2515_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2515_2 ( .OUT(na2515_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2515_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2515_4 ( .OUT(na2515_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2517_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2515_5 ( .OUT(na2515_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2515_2_i) );
// C_AND/D//AND/D      x20y38     80'h00_F600_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2517_1 ( .OUT(na2517_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2517_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2517_2 ( .OUT(na2517_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2517_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2517_4 ( .OUT(na2517_2_i), .IN1(1'b1), .IN2(na2519_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2517_5 ( .OUT(na2517_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2517_2_i) );
// C_AND/D//AND/D      x19y40     80'h00_F600_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2519_1 ( .OUT(na2519_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2519_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2519_2 ( .OUT(na2519_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2519_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2519_4 ( .OUT(na2519_2_i), .IN1(na2521_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2519_5 ( .OUT(na2519_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2519_2_i) );
// C_AND/D//AND/D      x17y39     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2521_1 ( .OUT(na2521_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2521_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2521_2 ( .OUT(na2521_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2521_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2521_4 ( .OUT(na2521_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2523_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2521_5 ( .OUT(na2521_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2521_2_i) );
// C_AND/D//AND/D      x18y41     80'h00_F600_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2523_1 ( .OUT(na2523_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2523_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2523_2 ( .OUT(na2523_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2523_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2523_4 ( .OUT(na2523_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2525_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2523_5 ( .OUT(na2523_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2523_2_i) );
// C_AND/D//AND/D      x16y44     80'h00_F600_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2525_1 ( .OUT(na2525_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2525_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2525_2 ( .OUT(na2525_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2525_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2525_4 ( .OUT(na2525_2_i), .IN1(1'b1), .IN2(na2527_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2525_5 ( .OUT(na2525_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2525_2_i) );
// C_AND/D//AND/D      x19y44     80'h00_F600_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2527_1 ( .OUT(na2527_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2527_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2527_2 ( .OUT(na2527_1), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2527_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2527_4 ( .OUT(na2527_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2529_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2527_5 ( .OUT(na2527_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2527_2_i) );
// C_///AND/D      x22y55     80'h00_F600_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2529_4 ( .OUT(na2529_2_i), .IN1(na886_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2529_5 ( .OUT(na2529_2), .CLK(na1739_1), .EN(~na1475_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2529_2_i) );
// C_AND/D//AND/D      x16y45     80'h00_FA00_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2579_1 ( .OUT(na2579_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2579_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2579_2 ( .OUT(na2579_1), .CLK(na1739_1), .EN(na1479_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2579_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2579_4 ( .OUT(na2579_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2581_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2579_5 ( .OUT(na2579_2), .CLK(na1739_1), .EN(na1479_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2579_2_i) );
// C_AND/D///      x16y48     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2581_1 ( .OUT(na2581_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na891_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2581_2 ( .OUT(na2581_1), .CLK(na1739_1), .EN(na1479_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2581_1_i) );
// C_AND/D//AND/D      x40y35     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2593_1 ( .OUT(na2593_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3531_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2593_2 ( .OUT(na2593_1), .CLK(na1739_1), .EN(na1415_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2593_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2593_4 ( .OUT(na2593_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3532_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2593_5 ( .OUT(na2593_2), .CLK(na1739_1), .EN(na1415_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2593_2_i) );
// C_AND/D//AND/D      x36y43     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2595_1 ( .OUT(na2595_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3529_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2595_2 ( .OUT(na2595_1), .CLK(na1739_1), .EN(na1415_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2595_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2595_4 ( .OUT(na2595_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3530_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2595_5 ( .OUT(na2595_2), .CLK(na1739_1), .EN(na1415_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2595_2_i) );
// C_AND/D//AND/D      x42y43     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2597_1 ( .OUT(na2597_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3527_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2597_2 ( .OUT(na2597_1), .CLK(na1739_1), .EN(na1415_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2597_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2597_4 ( .OUT(na2597_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3528_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2597_5 ( .OUT(na2597_2), .CLK(na1739_1), .EN(na1415_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2597_2_i) );
// C_AND/D//AND/D      x30y43     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2599_1 ( .OUT(na2599_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3525_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2599_2 ( .OUT(na2599_1), .CLK(na1739_1), .EN(na1415_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2599_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2599_4 ( .OUT(na2599_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3526_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2599_5 ( .OUT(na2599_2), .CLK(na1739_1), .EN(na1415_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2599_2_i) );
// C_AND/D//AND/D      x39y49     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2600_1 ( .OUT(na2600_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2600_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2600_2 ( .OUT(na2600_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2600_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2600_4 ( .OUT(na2600_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2602_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2600_5 ( .OUT(na2600_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2600_2_i) );
// C_AND/D//AND/D      x36y50     80'h00_FE00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2602_1 ( .OUT(na2602_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2602_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2602_2 ( .OUT(na2602_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2602_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2602_4 ( .OUT(na2602_2_i), .IN1(1'b1), .IN2(na2604_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2602_5 ( .OUT(na2602_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2602_2_i) );
// C_AND/D//AND/D      x31y50     80'h00_FE00_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2604_1 ( .OUT(na2604_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2604_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2604_2 ( .OUT(na2604_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2604_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2604_4 ( .OUT(na2604_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na951_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2604_5 ( .OUT(na2604_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2604_2_i) );
// C_///AND/D      x36y65     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2705_4 ( .OUT(na2705_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3414_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2705_5 ( .OUT(na2705_2), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2705_2_i) );
// C_AND/D///      x45y90     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2706_1 ( .OUT(na2706_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1784_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2706_2 ( .OUT(na2706_1), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2706_1_i) );
// C_AND/D//AND/D      x48y90     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2707_1 ( .OUT(na2707_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1784_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2707_2 ( .OUT(na2707_1), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2707_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2707_4 ( .OUT(na2707_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1786_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2707_5 ( .OUT(na2707_2), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2707_2_i) );
// C_///AND/D      x46y86     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2710_4 ( .OUT(na2710_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2842_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2710_5 ( .OUT(na2710_2), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2710_2_i) );
// C_AND/D//AND/D      x37y79     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2712_1 ( .OUT(na2712_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2844_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2712_2 ( .OUT(na2712_1), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2712_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2712_4 ( .OUT(na2712_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2844_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2712_5 ( .OUT(na2712_2), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2712_2_i) );
// C_AND/D//AND/D      x38y83     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2713_1 ( .OUT(na2713_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2846_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2713_2 ( .OUT(na2713_1), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2713_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2713_4 ( .OUT(na2713_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2842_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2713_5 ( .OUT(na2713_2), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2713_2_i) );
// C_AND/D///      x39y73     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2714_1 ( .OUT(na2714_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3413_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2714_2 ( .OUT(na2714_1), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2714_1_i) );
// C_///AND/D      x58y66     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2715_4 ( .OUT(na2715_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1792_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2715_5 ( .OUT(na2715_2), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2715_2_i) );
// C_AND/D///      x45y71     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2716_1 ( .OUT(na2716_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1792_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2716_2 ( .OUT(na2716_1), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2716_1_i) );
// C_///AND/D      x62y68     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2717_4 ( .OUT(na2717_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1794_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2717_5 ( .OUT(na2717_2), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2717_2_i) );
// C_AND/D///      x50y72     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2718_1 ( .OUT(na2718_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1794_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2718_2 ( .OUT(na2718_1), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2718_1_i) );
// C_///AND/D      x46y52     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2719_4 ( .OUT(na2719_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3424_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2719_5 ( .OUT(na2719_2), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2719_2_i) );
// C_AND/D///      x40y70     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2720_1 ( .OUT(na2720_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2846_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2720_2 ( .OUT(na2720_1), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2720_1_i) );
// C_///AND/D      x42y74     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2721_4 ( .OUT(na2721_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1780_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2721_5 ( .OUT(na2721_2), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2721_2_i) );
// C_AND/D//AND/D      x40y68     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2722_1 ( .OUT(na2722_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1780_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2722_2 ( .OUT(na2722_1), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2722_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2722_4 ( .OUT(na2722_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1782_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2722_5 ( .OUT(na2722_2), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2722_2_i) );
// C_///AND/D      x50y72     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2723_4 ( .OUT(na2723_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1782_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2723_5 ( .OUT(na2723_2), .CLK(na1739_1), .EN(na218_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2723_2_i) );
// C_///AND/D      x60y86     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2730_4 ( .OUT(na2730_2_i), .IN1(1'b1), .IN2(na1044_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2730_5 ( .OUT(na2730_2), .CLK(na1739_1), .EN(na1502_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2730_2_i) );
// C_AND/D//AND/D      x38y90     80'h00_F600_80_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2739_1 ( .OUT(na2739_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2739_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2739_2 ( .OUT(na2739_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2739_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2739_4 ( .OUT(na2739_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2741_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2739_5 ( .OUT(na2739_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2739_2_i) );
// C_AND/D//AND/D      x32y79     80'h00_F600_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2741_1 ( .OUT(na2741_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2741_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2741_2 ( .OUT(na2741_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2741_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2741_4 ( .OUT(na2741_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2743_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2741_5 ( .OUT(na2741_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2741_2_i) );
// C_AND/D//AND/D      x30y75     80'h00_F600_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2743_1 ( .OUT(na2743_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2743_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2743_2 ( .OUT(na2743_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2743_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2743_4 ( .OUT(na2743_2_i), .IN1(1'b1), .IN2(na2745_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2743_5 ( .OUT(na2743_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2743_2_i) );
// C_AND/D//AND/D      x21y74     80'h00_F600_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2745_1 ( .OUT(na2745_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2745_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2745_2 ( .OUT(na2745_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2745_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2745_4 ( .OUT(na2745_2_i), .IN1(na2747_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2745_5 ( .OUT(na2745_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2745_2_i) );
// C_AND/D//AND/D      x15y81     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2747_1 ( .OUT(na2747_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2747_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2747_2 ( .OUT(na2747_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2747_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2747_4 ( .OUT(na2747_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2749_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2747_5 ( .OUT(na2747_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2747_2_i) );
// C_AND/D//AND/D      x14y85     80'h00_F600_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2749_1 ( .OUT(na2749_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2749_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2749_2 ( .OUT(na2749_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2749_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2749_4 ( .OUT(na2749_2_i), .IN1(1'b1), .IN2(na2751_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2749_5 ( .OUT(na2749_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2749_2_i) );
// C_AND/D//AND/D      x15y88     80'h00_F600_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2751_1 ( .OUT(na2751_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2751_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2751_2 ( .OUT(na2751_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2751_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2751_4 ( .OUT(na2751_2_i), .IN1(1'b1), .IN2(na2753_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2751_5 ( .OUT(na2751_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2751_2_i) );
// C_AND/D//AND/D      x13y88     80'h00_F600_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2753_1 ( .OUT(na2753_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2753_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2753_2 ( .OUT(na2753_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2753_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2753_4 ( .OUT(na2753_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2755_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2753_5 ( .OUT(na2753_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2753_2_i) );
// C_AND/D//AND/D      x14y89     80'h00_F600_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2755_1 ( .OUT(na2755_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2755_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2755_2 ( .OUT(na2755_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2755_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2755_4 ( .OUT(na2755_2_i), .IN1(na2757_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2755_5 ( .OUT(na2755_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2755_2_i) );
// C_AND/D//AND/D      x15y89     80'h00_F600_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2757_1 ( .OUT(na2757_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2757_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2757_2 ( .OUT(na2757_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2757_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2757_4 ( .OUT(na2757_2_i), .IN1(1'b1), .IN2(na2759_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2757_5 ( .OUT(na2757_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2757_2_i) );
// C_AND/D//AND/D      x15y90     80'h00_F600_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2759_1 ( .OUT(na2759_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2759_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2759_2 ( .OUT(na2759_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2759_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2759_4 ( .OUT(na2759_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2761_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2759_5 ( .OUT(na2759_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2759_2_i) );
// C_AND/D//AND/D      x14y91     80'h00_F600_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2761_1 ( .OUT(na2761_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2761_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2761_2 ( .OUT(na2761_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2761_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2761_4 ( .OUT(na2761_2_i), .IN1(na2763_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2761_5 ( .OUT(na2761_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2761_2_i) );
// C_AND/D//AND/D      x15y91     80'h00_F600_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2763_1 ( .OUT(na2763_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2763_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2763_2 ( .OUT(na2763_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2763_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2763_4 ( .OUT(na2763_2_i), .IN1(1'b1), .IN2(na2765_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2763_5 ( .OUT(na2763_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2763_2_i) );
// C_AND/D//AND/D      x19y92     80'h00_F600_80_0000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2765_1 ( .OUT(na2765_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2765_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2765_2 ( .OUT(na2765_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2765_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2765_4 ( .OUT(na2765_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2767_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2765_5 ( .OUT(na2765_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2765_2_i) );
// C_AND/D//AND/D      x32y91     80'h00_F600_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2767_1 ( .OUT(na2767_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2767_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2767_2 ( .OUT(na2767_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2767_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2767_4 ( .OUT(na2767_2_i), .IN1(na2769_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2767_5 ( .OUT(na2767_2), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2767_2_i) );
// C_AND/D///      x47y87     80'h00_F600_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2769_1 ( .OUT(na2769_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1050_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2769_2 ( .OUT(na2769_1), .CLK(na1739_1), .EN(~na1497_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2769_1_i) );
// C_AND/D//AND/D      x19y91     80'h00_FA00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2819_1 ( .OUT(na2819_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2819_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2819_2 ( .OUT(na2819_1), .CLK(na1739_1), .EN(na1501_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2819_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2819_4 ( .OUT(na2819_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2821_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2819_5 ( .OUT(na2819_2), .CLK(na1739_1), .EN(na1501_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2819_2_i) );
// C_///AND/D      x22y92     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2821_4 ( .OUT(na2821_2_i), .IN1(1'b1), .IN2(na1051_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2821_5 ( .OUT(na2821_2), .CLK(na1739_1), .EN(na1501_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2821_2_i) );
// C_AND/D//AND/D      x46y56     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2840_1 ( .OUT(na2840_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3423_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2840_2 ( .OUT(na2840_1), .CLK(na1739_1), .EN(na1419_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2840_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2840_4 ( .OUT(na2840_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3424_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2840_5 ( .OUT(na2840_2), .CLK(na1739_1), .EN(na1419_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2840_2_i) );
// C_AND/D//AND/D      x46y68     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2842_1 ( .OUT(na2842_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3420_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2842_2 ( .OUT(na2842_1), .CLK(na1739_1), .EN(na1419_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2842_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2842_4 ( .OUT(na2842_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3421_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2842_5 ( .OUT(na2842_2), .CLK(na1739_1), .EN(na1419_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2842_2_i) );
// C_AND/D//AND/D      x44y68     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2844_1 ( .OUT(na2844_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3416_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2844_2 ( .OUT(na2844_1), .CLK(na1739_1), .EN(na1419_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2844_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2844_4 ( .OUT(na2844_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3417_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2844_5 ( .OUT(na2844_2), .CLK(na1739_1), .EN(na1419_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2844_2_i) );
// C_AND/D//AND/D      x44y70     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2846_1 ( .OUT(na2846_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3413_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2846_2 ( .OUT(na2846_1), .CLK(na1739_1), .EN(na1419_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2846_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2846_4 ( .OUT(na2846_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3414_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2846_5 ( .OUT(na2846_2), .CLK(na1739_1), .EN(na1419_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2846_2_i) );
// C_AND/D//AND/D      x60y91     80'h00_FE00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2847_1 ( .OUT(na2847_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2847_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2847_2 ( .OUT(na2847_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2847_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2847_4 ( .OUT(na2847_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2849_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2847_5 ( .OUT(na2847_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2847_2_i) );
// C_AND/D//AND/D      x60y89     80'h00_FE00_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2849_1 ( .OUT(na2849_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2849_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2849_2 ( .OUT(na2849_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2849_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2849_4 ( .OUT(na2849_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2851_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2849_5 ( .OUT(na2849_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2849_2_i) );
// C_AND/D//AND/D      x54y90     80'h00_FE00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2851_1 ( .OUT(na2851_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2851_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2851_2 ( .OUT(na2851_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2851_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2851_4 ( .OUT(na2851_2_i), .IN1(1'b1), .IN2(na1112_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2851_5 ( .OUT(na2851_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na2851_2_i) );
// C_AND/D///      x49y63     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2956_1 ( .OUT(na2956_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3427_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2956_2 ( .OUT(na2956_1), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2956_1_i) );
// C_///AND/D      x65y87     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2957_4 ( .OUT(na2957_2_i), .IN1(1'b1), .IN2(na1767_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2957_5 ( .OUT(na2957_2), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2957_2_i) );
// C_AND/D//AND/D      x62y85     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2958_1 ( .OUT(na2958_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1767_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2958_2 ( .OUT(na2958_1), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2958_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2958_4 ( .OUT(na2958_2_i), .IN1(1'b1), .IN2(na1769_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2958_5 ( .OUT(na2958_2), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2958_2_i) );
// C_AND/D///      x62y83     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2961_1 ( .OUT(na2961_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3100_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2961_2 ( .OUT(na2961_1), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2961_1_i) );
// C_AND/D//AND/D      x55y83     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2962_1 ( .OUT(na2962_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3102_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2962_2 ( .OUT(na2962_1), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2962_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2962_4 ( .OUT(na2962_2_i), .IN1(1'b1), .IN2(na3100_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2962_5 ( .OUT(na2962_2), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2962_2_i) );
// C_///AND/D      x59y83     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2963_4 ( .OUT(na2963_2_i), .IN1(1'b1), .IN2(na3102_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2963_5 ( .OUT(na2963_2), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2963_2_i) );
// C_AND/D//AND/D      x51y82     80'h00_FA00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2965_1 ( .OUT(na2965_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3426_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2965_2 ( .OUT(na2965_1), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2965_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2965_4 ( .OUT(na2965_2_i), .IN1(1'b1), .IN2(na3104_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2965_5 ( .OUT(na2965_2), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2965_2_i) );
// C_AND/D///      x33y58     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2966_1 ( .OUT(na2966_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1775_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2966_2 ( .OUT(na2966_1), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2966_1_i) );
// C_///AND/D      x33y54     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2967_4 ( .OUT(na2967_2_i), .IN1(1'b1), .IN2(na1775_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2967_5 ( .OUT(na2967_2), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2967_2_i) );
// C_AND/D///      x34y57     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2968_1 ( .OUT(na2968_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1777_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2968_2 ( .OUT(na2968_1), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2968_1_i) );
// C_///AND/D      x33y49     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2969_4 ( .OUT(na2969_2_i), .IN1(1'b1), .IN2(na1777_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2969_5 ( .OUT(na2969_2), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2969_2_i) );
// C_AND/D///      x30y46     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2970_1 ( .OUT(na2970_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3444_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2970_2 ( .OUT(na2970_1), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2970_1_i) );
// C_///AND/D      x32y58     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2971_4 ( .OUT(na2971_2_i), .IN1(1'b1), .IN2(na3104_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2971_5 ( .OUT(na2971_2), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2971_2_i) );
// C_AND/D///      x28y63     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2972_1 ( .OUT(na2972_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1763_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2972_2 ( .OUT(na2972_1), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2972_1_i) );
// C_AND/D//AND/D      x25y62     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2973_1 ( .OUT(na2973_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1763_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2973_2 ( .OUT(na2973_1), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2973_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2973_4 ( .OUT(na2973_2_i), .IN1(1'b1), .IN2(na1765_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2973_5 ( .OUT(na2973_2), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2973_2_i) );
// C_///AND/D      x29y63     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2974_4 ( .OUT(na2974_2_i), .IN1(1'b1), .IN2(na1765_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2974_5 ( .OUT(na2974_2), .CLK(na1739_1), .EN(na436_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2974_2_i) );
// C_AND/D///      x57y84     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2981_1 ( .OUT(na2981_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1192_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2981_2 ( .OUT(na2981_1), .CLK(na1739_1), .EN(na1524_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2981_1_i) );
// C_AND/D//AND/D      x48y87     80'h00_F600_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2984_1 ( .OUT(na2984_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2984_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2984_2 ( .OUT(na2984_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2984_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2984_4 ( .OUT(na2984_2_i), .IN1(na2986_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2984_5 ( .OUT(na2984_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2984_2_i) );
// C_AND/D//AND/D      x23y71     80'h00_F600_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2986_1 ( .OUT(na2986_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2986_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2986_2 ( .OUT(na2986_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2986_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2986_4 ( .OUT(na2986_2_i), .IN1(na2988_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2986_5 ( .OUT(na2986_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2986_2_i) );
// C_AND/D//AND/D      x15y73     80'h00_F600_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2988_1 ( .OUT(na2988_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2988_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2988_2 ( .OUT(na2988_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2988_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2988_4 ( .OUT(na2988_2_i), .IN1(1'b1), .IN2(na2990_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2988_5 ( .OUT(na2988_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2988_2_i) );
// C_AND/D//AND/D      x13y74     80'h00_F600_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2990_1 ( .OUT(na2990_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2990_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2990_2 ( .OUT(na2990_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2990_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2990_4 ( .OUT(na2990_2_i), .IN1(na2992_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2990_5 ( .OUT(na2990_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2990_2_i) );
// C_AND/D//AND/D      x13y79     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2992_1 ( .OUT(na2992_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2992_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2992_2 ( .OUT(na2992_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2992_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2992_4 ( .OUT(na2992_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na2994_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2992_5 ( .OUT(na2992_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2992_2_i) );
// C_AND/D//AND/D      x14y81     80'h00_F600_80_0000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2994_1 ( .OUT(na2994_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2994_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2994_2 ( .OUT(na2994_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2994_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2994_4 ( .OUT(na2994_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na2996_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2994_5 ( .OUT(na2994_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2994_2_i) );
// C_AND/D//AND/D      x14y78     80'h00_F600_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2996_1 ( .OUT(na2996_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na2996_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2996_2 ( .OUT(na2996_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2996_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2996_4 ( .OUT(na2996_2_i), .IN1(na2998_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2996_5 ( .OUT(na2996_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2996_2_i) );
// C_AND/D//AND/D      x15y75     80'h00_F600_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a2998_1 ( .OUT(na2998_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2998_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a2998_2 ( .OUT(na2998_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2998_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a2998_4 ( .OUT(na2998_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3000_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a2998_5 ( .OUT(na2998_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na2998_2_i) );
// C_AND/D//AND/D      x14y71     80'h00_F600_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3000_1 ( .OUT(na3000_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3000_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3000_2 ( .OUT(na3000_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3000_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3000_4 ( .OUT(na3000_2_i), .IN1(na3002_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3000_5 ( .OUT(na3000_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3000_2_i) );
// C_AND/D//AND/D      x15y69     80'h00_F600_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3002_1 ( .OUT(na3002_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3002_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3002_2 ( .OUT(na3002_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3002_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3002_4 ( .OUT(na3002_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3004_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3002_5 ( .OUT(na3002_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3002_2_i) );
// C_AND/D//AND/D      x14y70     80'h00_F600_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3004_1 ( .OUT(na3004_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3004_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3004_2 ( .OUT(na3004_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3004_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3004_4 ( .OUT(na3004_2_i), .IN1(na3006_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3004_5 ( .OUT(na3004_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3004_2_i) );
// C_AND/D//AND/D      x13y75     80'h00_F600_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3006_1 ( .OUT(na3006_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3006_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3006_2 ( .OUT(na3006_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3006_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3006_4 ( .OUT(na3006_2_i), .IN1(1'b1), .IN2(na3008_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3006_5 ( .OUT(na3006_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3006_2_i) );
// C_AND/D//AND/D      x15y78     80'h00_F600_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3008_1 ( .OUT(na3008_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na3008_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3008_2 ( .OUT(na3008_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3008_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3008_4 ( .OUT(na3008_2_i), .IN1(na3010_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3008_5 ( .OUT(na3008_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3008_2_i) );
// C_AND/D//AND/D      x15y79     80'h00_F600_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3010_1 ( .OUT(na3010_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3010_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3010_2 ( .OUT(na3010_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3010_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3010_4 ( .OUT(na3010_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3012_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3010_5 ( .OUT(na3010_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3010_2_i) );
// C_AND/D//AND/D      x22y76     80'h00_F600_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3012_1 ( .OUT(na3012_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3012_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3012_2 ( .OUT(na3012_1), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3012_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3012_4 ( .OUT(na3012_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3014_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3012_5 ( .OUT(na3012_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3012_2_i) );
// C_///AND/D      x44y76     80'h00_F600_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3014_4 ( .OUT(na3014_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1198_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3014_5 ( .OUT(na3014_2), .CLK(na1739_1), .EN(~na1519_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3014_2_i) );
// C_AND/D//AND/D      x70y91     80'h00_FA00_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3064_1 ( .OUT(na3064_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3064_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3064_2 ( .OUT(na3064_1), .CLK(na1739_1), .EN(na1523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3064_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3064_4 ( .OUT(na3064_2_i), .IN1(1'b1), .IN2(na3066_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3064_5 ( .OUT(na3064_2), .CLK(na1739_1), .EN(na1523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3064_2_i) );
// C_AND/D///      x67y92     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3066_1 ( .OUT(na3066_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1199_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3066_2 ( .OUT(na3066_1), .CLK(na1739_1), .EN(na1523_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3066_1_i) );
// C_AND/D//AND/D      x37y50     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3098_1 ( .OUT(na3098_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3443_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3098_2 ( .OUT(na3098_1), .CLK(na1739_1), .EN(na1422_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3098_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3098_4 ( .OUT(na3098_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3444_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3098_5 ( .OUT(na3098_2), .CLK(na1739_1), .EN(na1422_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3098_2_i) );
// C_AND/D//AND/D      x43y58     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3100_1 ( .OUT(na3100_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3439_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3100_2 ( .OUT(na3100_1), .CLK(na1739_1), .EN(na1422_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3100_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3100_4 ( .OUT(na3100_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3442_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3100_5 ( .OUT(na3100_2), .CLK(na1739_1), .EN(na1422_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3100_2_i) );
// C_AND/D//AND/D      x41y56     80'h00_FA00_80_0000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3102_1 ( .OUT(na3102_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na3429_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3102_2 ( .OUT(na3102_1), .CLK(na1739_1), .EN(na1422_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3102_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3102_4 ( .OUT(na3102_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na3430_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3102_5 ( .OUT(na3102_2), .CLK(na1739_1), .EN(na1422_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3102_2_i) );
// C_AND/D//AND/D      x43y56     80'h00_FA00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3104_1 ( .OUT(na3104_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3426_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3104_2 ( .OUT(na3104_1), .CLK(na1739_1), .EN(na1422_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3104_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3104_4 ( .OUT(na3104_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3427_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3104_5 ( .OUT(na3104_2), .CLK(na1739_1), .EN(na1422_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0),
                      .D_IN(na3104_2_i) );
// C_AND/D//AND/D      x43y63     80'h00_FE00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3105_1 ( .OUT(na3105_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3105_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3105_2 ( .OUT(na3105_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3105_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3105_4 ( .OUT(na3105_2_i), .IN1(na3107_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3105_5 ( .OUT(na3105_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3105_2_i) );
// C_AND/D//AND/D      x43y65     80'h00_FE00_80_0000_0C88_FACF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3107_1 ( .OUT(na3107_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3107_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3107_2 ( .OUT(na3107_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3107_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3107_4 ( .OUT(na3107_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na3109_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3107_5 ( .OUT(na3107_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3107_2_i) );
// C_AND/D//AND/D      x46y72     80'h00_FE00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3109_1 ( .OUT(na3109_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na3109_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a3109_2 ( .OUT(na3109_1), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3109_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3109_4 ( .OUT(na3109_2_i), .IN1(1'b1), .IN2(na1254_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a3109_5 ( .OUT(na3109_2), .CLK(na1739_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na3109_2_i) );
// C_MX4b////      x51y77     80'h00_0018_00_0040_0AFE_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3145_1 ( .OUT(na3145_1), .IN1(1'b1), .IN2(na1541_2), .IN3(na4461_2), .IN4(1'b1), .IN5(na1429_2), .IN6(~na1536_1), .IN7(~na1537_2),
                      .IN8(~na1538_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x52y87     80'h00_0018_00_0040_0AFD_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3146_1 ( .OUT(na3146_1), .IN1(1'b1), .IN2(~na1543_2), .IN3(na4465_2), .IN4(1'b1), .IN5(~na1514_2), .IN6(na1428_1), .IN7(~na1516_2),
                      .IN8(~na1515_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x13y68     80'h00_0018_00_0040_0A55_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3147_1 ( .OUT(na3147_1), .IN1(1'b1), .IN2(na24_1), .IN3(~na233_2), .IN4(1'b1), .IN5(~na1614_2), .IN6(1'b0), .IN7(~na4472_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x17y68     80'h00_0018_00_0040_0AA0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3148_1 ( .OUT(na3148_1), .IN1(1'b1), .IN2(~na24_1), .IN3(~na233_2), .IN4(1'b1), .IN5(1'b0), .IN6(na155_2), .IN7(1'b0), .IN8(na156_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x17y69     80'h00_0018_00_0040_0A50_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3149_1 ( .OUT(na3149_1), .IN1(1'b1), .IN2(na24_1), .IN3(na233_2), .IN4(1'b1), .IN5(na235_2), .IN6(1'b0), .IN7(na233_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x16y70     80'h00_0018_00_0040_0A50_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3150_1 ( .OUT(na3150_1), .IN1(1'b1), .IN2(na24_1), .IN3(~na233_2), .IN4(1'b1), .IN5(na234_1), .IN6(1'b0), .IN7(na236_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y59     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3151_1 ( .OUT(na3151_1), .IN1(na1314_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4154_2), .IN5(na1200_1), .IN6(na1052_1), .IN7(na892_1),
                      .IN8(na728_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y55     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3152_1 ( .OUT(na3152_1), .IN1(na1314_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4154_2), .IN5(na1200_2), .IN6(na1052_2), .IN7(na892_2),
                      .IN8(na728_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y60     80'h00_0018_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3153_1 ( .OUT(na3153_1), .IN1(~na1314_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4154_2), .IN5(na1054_1), .IN6(na4375_2), .IN7(na730_1),
                      .IN8(na4306_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x49y60     80'h00_0018_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3154_1 ( .OUT(na3154_1), .IN1(~na1314_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4154_2), .IN5(na1054_2), .IN6(na4376_2), .IN7(na730_2),
                      .IN8(na4307_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y65     80'h00_0018_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3155_1 ( .OUT(na3155_1), .IN1(~na1314_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4154_2), .IN5(na1056_1), .IN6(na1204_1), .IN7(na732_1),
                      .IN8(na896_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x52y62     80'h00_0018_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3156_1 ( .OUT(na3156_1), .IN1(~na1314_2), .IN2(1'b1), .IN3(1'b1), .IN4(na4154_2), .IN5(na1056_2), .IN6(na1204_2), .IN7(na732_2),
                      .IN8(na896_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y60     80'h00_0018_00_0040_0AF0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3157_1 ( .OUT(na3157_1), .IN1(~na1314_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4154_2), .IN5(na734_1), .IN6(na898_1), .IN7(na1058_1),
                      .IN8(na1206_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y64     80'h00_0018_00_0040_0AF0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3158_1 ( .OUT(na3158_1), .IN1(~na1314_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4154_2), .IN5(na734_2), .IN6(na898_2), .IN7(na1058_2),
                      .IN8(na1206_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x49y72     80'h00_0018_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3159_1 ( .OUT(na3159_1), .IN1(na1314_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4154_2), .IN5(na4067_2), .IN6(na4_1), .IN7(na8_1),
                      .IN8(na4066_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x18y67     80'h00_0018_00_0040_0A55_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3160_1 ( .OUT(na3160_1), .IN1(1'b1), .IN2(na24_1), .IN3(~na233_2), .IN4(1'b1), .IN5(~na394_1), .IN6(1'b0), .IN7(~na395_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x18y73     80'h00_0018_00_0040_0A50_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3161_1 ( .OUT(na3161_1), .IN1(1'b1), .IN2(~na25_2), .IN3(~na233_2), .IN4(1'b1), .IN5(na1148_2), .IN6(1'b0), .IN7(na1316_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x70y44     80'h00_0018_00_0040_0AFE_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3162_1 ( .OUT(na3162_1), .IN1(1'b1), .IN2(na1542_2), .IN3(1'b1), .IN4(na4463_2), .IN5(na1426_2), .IN6(~na1470_1), .IN7(~na1471_2),
                      .IN8(~na1472_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x66y65     80'h00_0060_00_0000_0C06_FFC9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3163_4 ( .OUT(na3163_2), .IN1(na535_1), .IN2(~na512_1), .IN3(1'b0), .IN4(na1985_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x65y67     80'h00_0018_00_0040_0A67_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3164_1 ( .OUT(na3164_1), .IN1(~na535_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1985_1), .IN5(1'b1), .IN6(~na512_1), .IN7(~na4215_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x67y48     80'h00_0018_00_0040_0AF0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3165_1 ( .OUT(na3165_1), .IN1(~na4467_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1544_1), .IN5(na567_1), .IN6(na559_1), .IN7(na551_1),
                      .IN8(na4229_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x69y48     80'h00_0018_00_0040_0AF0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3166_1 ( .OUT(na3166_1), .IN1(~na4467_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1544_1), .IN5(na567_2), .IN6(na559_2), .IN7(na551_2),
                      .IN8(na4230_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x63y45     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3167_1 ( .OUT(na3167_1), .IN1(na4467_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1544_1), .IN5(na545_1), .IN6(na553_1), .IN7(na561_1),
                      .IN8(na4247_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x65y46     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3168_1 ( .OUT(na3168_1), .IN1(na4467_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1544_1), .IN5(na545_2), .IN6(na553_2), .IN7(na561_2),
                      .IN8(na4248_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x66y45     80'h00_0018_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3169_1 ( .OUT(na3169_1), .IN1(na4467_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1544_1), .IN5(na563_1), .IN6(na4249_2), .IN7(na547_1),
                      .IN8(na4239_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x70y46     80'h00_0018_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3170_1 ( .OUT(na3170_1), .IN1(na4467_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1544_1), .IN5(na563_2), .IN6(na4250_2), .IN7(na547_2),
                      .IN8(na4240_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x64y46     80'h00_0018_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3171_1 ( .OUT(na3171_1), .IN1(na4467_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1544_1), .IN5(na565_1), .IN6(na4251_2), .IN7(na549_1),
                      .IN8(na4241_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x63y46     80'h00_0018_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3172_1 ( .OUT(na3172_1), .IN1(na4467_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1544_1), .IN5(na565_2), .IN6(na4252_2), .IN7(na549_2),
                      .IN8(na4242_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x20y74     80'h00_0018_00_0040_0C05_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3173_1 ( .OUT(na3173_1), .IN1(na643_2), .IN2(1'b0), .IN3(na644_1), .IN4(1'b0), .IN5(1'b1), .IN6(na25_2), .IN7(~na233_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x18y74     80'h00_0018_00_0040_0C0A_5300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3174_1 ( .OUT(na3174_1), .IN1(1'b0), .IN2(na687_2), .IN3(1'b0), .IN4(na689_1), .IN5(1'b1), .IN6(~na25_2), .IN7(~na233_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x63y51     80'h00_0018_00_0000_0C66_9A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3175_1 ( .OUT(na3175_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2222_1), .IN6(1'b0), .IN7(~na353_1), .IN8(na720_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x62y51     80'h00_0018_00_0040_0A67_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3176_1 ( .OUT(na3176_1), .IN1(na2222_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na720_1), .IN5(1'b1), .IN6(~na4175_2), .IN7(~na353_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x66y37     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3177_1 ( .OUT(na3177_1), .IN1(1'b1), .IN2(~na1542_2), .IN3(1'b1), .IN4(~na4463_2), .IN5(na752_1), .IN6(na4277_2), .IN7(na736_1),
                      .IN8(na728_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x64y38     80'h00_0018_00_0040_0AF0_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3178_1 ( .OUT(na3178_1), .IN1(1'b1), .IN2(~na1542_2), .IN3(1'b1), .IN4(~na4463_2), .IN5(na752_2), .IN6(na4278_2), .IN7(na736_2),
                      .IN8(na728_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x64y37     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3179_1 ( .OUT(na3179_1), .IN1(1'b1), .IN2(na1542_2), .IN3(1'b1), .IN4(~na4463_2), .IN5(na4279_2), .IN6(na754_1), .IN7(na730_1),
                      .IN8(na4271_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x66y38     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3180_1 ( .OUT(na3180_1), .IN1(1'b1), .IN2(na1542_2), .IN3(1'b1), .IN4(~na4463_2), .IN5(na4280_2), .IN6(na754_2), .IN7(na730_2),
                      .IN8(na4272_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x65y39     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3181_1 ( .OUT(na3181_1), .IN1(1'b1), .IN2(na1542_2), .IN3(1'b1), .IN4(~na4463_2), .IN5(na4281_2), .IN6(na756_1), .IN7(na732_1),
                      .IN8(na4273_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x66y40     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3182_1 ( .OUT(na3182_1), .IN1(1'b1), .IN2(na1542_2), .IN3(1'b1), .IN4(~na4463_2), .IN5(na4282_2), .IN6(na756_2), .IN7(na732_2),
                      .IN8(na4274_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x64y39     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3183_1 ( .OUT(na3183_1), .IN1(1'b1), .IN2(na1542_2), .IN3(1'b1), .IN4(na4463_2), .IN5(na734_1), .IN6(na4275_2), .IN7(na750_1),
                      .IN8(na4289_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x63y40     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3184_1 ( .OUT(na3184_1), .IN1(1'b1), .IN2(na1542_2), .IN3(1'b1), .IN4(na4463_2), .IN5(na734_2), .IN6(na4276_2), .IN7(na750_2),
                      .IN8(na4290_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x26y53     80'h00_0018_00_0000_0C66_C900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3185_1 ( .OUT(na3185_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na4296_2), .IN6(~na878_1), .IN7(1'b0), .IN8(na2473_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x26y56     80'h00_0018_00_0040_0A67_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3186_1 ( .OUT(na3186_1), .IN1(na4520_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na864_1), .IN5(1'b1), .IN6(~na878_1), .IN7(~na4298_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x43y43     80'h00_0018_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3187_1 ( .OUT(na3187_1), .IN1(na4468_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1545_1), .IN5(na908_1), .IN6(na916_1), .IN7(na892_1),
                      .IN8(na4310_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y44     80'h00_0018_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3188_1 ( .OUT(na3188_1), .IN1(na4468_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1545_1), .IN5(na908_2), .IN6(na916_2), .IN7(na892_2),
                      .IN8(na4311_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x41y42     80'h00_0018_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3189_1 ( .OUT(na3189_1), .IN1(~na4468_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1545_1), .IN5(na4312_2), .IN6(na894_1), .IN7(na918_1),
                      .IN8(na4320_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x42y42     80'h00_0018_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3190_1 ( .OUT(na3190_1), .IN1(~na4468_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1545_1), .IN5(na4313_2), .IN6(na894_2), .IN7(na918_2),
                      .IN8(na4321_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x43y44     80'h00_0018_00_0040_0AF0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3191_1 ( .OUT(na3191_1), .IN1(~na4468_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1545_1), .IN5(na4326_2), .IN6(na912_1), .IN7(na4314_2),
                      .IN8(na896_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x39y44     80'h00_0018_00_0040_0AF0_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3192_1 ( .OUT(na3192_1), .IN1(~na4468_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1545_1), .IN5(na4327_2), .IN6(na912_2), .IN7(na4315_2),
                      .IN8(na896_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x35y46     80'h00_0018_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3193_1 ( .OUT(na3193_1), .IN1(~na4468_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1545_1), .IN5(na4316_2), .IN6(na898_1), .IN7(na922_1),
                      .IN8(na4322_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x43y52     80'h00_0018_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3194_1 ( .OUT(na3194_1), .IN1(~na4468_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1545_1), .IN5(na4317_2), .IN6(na898_2), .IN7(na922_2),
                      .IN8(na4323_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x23y69     80'h00_0018_00_0040_0C05_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3195_1 ( .OUT(na3195_1), .IN1(na983_2), .IN2(1'b0), .IN3(na982_2), .IN4(1'b0), .IN5(1'b1), .IN6(na25_2), .IN7(na233_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x69y62     80'h00_0018_00_0040_0AF7_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3196_1 ( .OUT(na3196_1), .IN1(~na4467_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1544_1), .IN5(~na1450_2), .IN6(~na1449_2), .IN7(~na1448_1),
                      .IN8(na1425_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x39y86     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3197_1 ( .OUT(na3197_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2706_1), .IN7(~na1038_1), .IN8(na993_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x36y84     80'h00_0018_00_0040_0A67_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3198_1 ( .OUT(na3198_1), .IN1(1'b1), .IN2(na2706_1), .IN3(1'b1), .IN4(~na993_1), .IN5(1'b1), .IN6(~na4338_2), .IN7(~na1038_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y75     80'h00_0018_00_0040_0AF0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3199_1 ( .OUT(na3199_1), .IN1(1'b1), .IN2(~na1543_2), .IN3(na4465_2), .IN4(1'b1), .IN5(na1060_1), .IN6(na1052_1), .IN7(na4357_2),
                      .IN8(na4351_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x56y73     80'h00_0018_00_0040_0AF0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3200_1 ( .OUT(na3200_1), .IN1(1'b1), .IN2(~na1543_2), .IN3(na4465_2), .IN4(1'b1), .IN5(na1060_2), .IN6(na1052_2), .IN7(na4358_2),
                      .IN8(na4352_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x56y76     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3201_1 ( .OUT(na3201_1), .IN1(1'b1), .IN2(na1543_2), .IN3(na4465_2), .IN4(1'b1), .IN5(na1054_1), .IN6(na4344_2), .IN7(na4353_2),
                      .IN8(na4359_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y74     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3202_1 ( .OUT(na3202_1), .IN1(1'b1), .IN2(na1543_2), .IN3(na4465_2), .IN4(1'b1), .IN5(na1054_2), .IN6(na4345_2), .IN7(na4354_2),
                      .IN8(na4360_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y78     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3203_1 ( .OUT(na3203_1), .IN1(1'b1), .IN2(na1543_2), .IN3(na4465_2), .IN4(1'b1), .IN5(na1056_1), .IN6(na4346_2), .IN7(na4355_2),
                      .IN8(na1080_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y78     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3204_1 ( .OUT(na3204_1), .IN1(1'b1), .IN2(na1543_2), .IN3(na4465_2), .IN4(1'b1), .IN5(na1056_2), .IN6(na4347_2), .IN7(na4356_2),
                      .IN8(na1080_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x54y76     80'h00_0018_00_0040_0AF0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3205_1 ( .OUT(na3205_1), .IN1(1'b1), .IN2(na1543_2), .IN3(~na4465_2), .IN4(1'b1), .IN5(na1074_1), .IN6(na4363_2), .IN7(na1058_1),
                      .IN8(na4348_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y75     80'h00_0018_00_0040_0AF0_005C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3206_1 ( .OUT(na3206_1), .IN1(1'b1), .IN2(na1543_2), .IN3(~na4465_2), .IN4(1'b1), .IN5(na1074_2), .IN6(na4364_2), .IN7(na1058_2),
                      .IN8(na4349_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x61y77     80'h00_0018_00_0000_0C66_9A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3207_1 ( .OUT(na3207_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2957_2), .IN6(1'b0), .IN7(~na461_1), .IN8(na1388_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x61y82     80'h00_0018_00_0040_0A67_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3208_1 ( .OUT(na3208_1), .IN1(na2957_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1388_1), .IN5(1'b1), .IN6(~na4209_2), .IN7(~na461_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x40y59     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3209_1 ( .OUT(na3209_1), .IN1(1'b1), .IN2(na1541_2), .IN3(na4461_2), .IN4(1'b1), .IN5(na1200_1), .IN6(na4379_2), .IN7(na4387_2),
                      .IN8(na1224_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x37y58     80'h00_0018_00_0040_0AF0_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3210_1 ( .OUT(na3210_1), .IN1(1'b1), .IN2(na1541_2), .IN3(na4461_2), .IN4(1'b1), .IN5(na1200_2), .IN6(na4380_2), .IN7(na4388_2),
                      .IN8(na1224_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x37y64     80'h00_0018_00_0040_0AF0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3211_1 ( .OUT(na3211_1), .IN1(1'b1), .IN2(~na1541_2), .IN3(na4461_2), .IN4(1'b1), .IN5(na1210_1), .IN6(na4375_2), .IN7(na1226_1),
                      .IN8(na1218_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x32y55     80'h00_0018_00_0040_0AF0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3212_1 ( .OUT(na3212_1), .IN1(1'b1), .IN2(~na1541_2), .IN3(na4461_2), .IN4(1'b1), .IN5(na1210_2), .IN6(na4376_2), .IN7(na1226_2),
                      .IN8(na1218_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x33y59     80'h00_0018_00_0040_0AF0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3213_1 ( .OUT(na3213_1), .IN1(1'b1), .IN2(~na1541_2), .IN3(na4461_2), .IN4(1'b1), .IN5(na4383_2), .IN6(na1204_1), .IN7(na4394_2),
                      .IN8(na1220_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x35y60     80'h00_0018_00_0040_0AF0_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3214_1 ( .OUT(na3214_1), .IN1(1'b1), .IN2(~na1541_2), .IN3(na4461_2), .IN4(1'b1), .IN5(na4384_2), .IN6(na1204_2), .IN7(na4395_2),
                      .IN8(na1220_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x35y64     80'h00_0018_00_0040_0AF0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3215_1 ( .OUT(na3215_1), .IN1(1'b1), .IN2(~na1541_2), .IN3(~na4461_2), .IN4(1'b1), .IN5(na1230_1), .IN6(na4389_2), .IN7(na4385_2),
                      .IN8(na1206_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x34y61     80'h00_0018_00_0040_0AF0_0053
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3216_1 ( .OUT(na3216_1), .IN1(1'b1), .IN2(~na1541_2), .IN3(~na4461_2), .IN4(1'b1), .IN5(na1230_2), .IN6(na4390_2), .IN7(na4386_2),
                      .IN8(na1206_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x17y74     80'h00_0018_00_0040_0C05_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3217_1 ( .OUT(na3217_1), .IN1(na1148_2), .IN2(1'b0), .IN3(na1316_1), .IN4(1'b0), .IN5(1'b1), .IN6(na25_2), .IN7(~na233_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x35y49     80'h00_0018_00_0040_0AFE_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3218_1 ( .OUT(na3218_1), .IN1(na4468_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1545_1), .IN5(na1427_2), .IN6(~na1492_1), .IN7(~na1493_2),
                      .IN8(~na1494_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a3219 ( .Y(na3219_1), .I(i_clk) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a3220 ( .Y(na3220_1), .I(i_rstn) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010902)) 
           _a3221 ( .O(o_uart_tx), .A(na4065_10) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_0A_08_08_20_82),
             .REF_CLK(10.00),
             .OUT_CLK(16.00),
             .LOW_JITTER(1),
             .CI_FILTER_CONST(0),
             .CP_FILTER_CONST(0)) 
           _a3222 ( .USR_PLL_LOCKED_STDY(_d6), .USR_PLL_LOCKED(na3222_2), .CLK270(na3222_3), .CLK180(na3222_4), .CLK90(na3222_5), .CLK0(na3222_6),
                    .CLK_REF_OUT(_d7), .CLK_REF(na3229_1), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_0F_04_80_00_91_03_13_23_03_13_23_00_13_23_00_13_23_00_00),
             .INIT_00(320'h30000014b730000014b700cc50141300cc5014130000001417000000141700000000130000000013),
             .INIT_01(320'h00015014130001501413000050088300005008830005520023000552002302c700089302c7000893),
             .INIT_02(320'h00000088b700000088b700055240230005524023040023889304002388933f802268e33f802268e3),
             .INIT_03(320'h3f05f3c06f3f05f3c06f3f802278e33f802278e33fcf2208933fcf2208931c402208931c40220893),
             .INIT_04(320'h080731e461080731e4611cc200c4301cc200c0300c0300c0200c0300c020194721bc43194721bc43),
             .INIT_05(320'h0000000000000000000000000000000000000000000000286f000000286f1b06c194681b06c19468),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a3223 ( .DOA({_d8, _d9, _d10, _d11, _d12, _d13, _d14, _d15, _d16, _d17, _d18, _d19, _d20, _d21, _d22, _d23, _d24, _d25,
                   _d26, _d27, _d28, _d29, _d30, _d31, _d32, _d33, _d34, _d35, _d36, _d37, _d38, _d39, _d40, _d41, _d42, _d43, _d44,
                   _d45, _d46, _d47}),
                    .DOAX({_d48, _d49, _d50, _d51, _d52, _d53, _d54, _d55, _d56, _d57, _d58, _d59, _d60, _d61, _d62, _d63, _d64, _d65,
                   _d66, _d67, _d68, _d69, _d70, _d71, _d72, _d73, _d74, _d75, _d76, _d77, _d78, _d79, _d80, _d81, _d82, _d83, _d84,
                   _d85, _d86, _d87}),
                    .DOB({_d88, _d89, _d90, _d91, _d92, _d93, _d94, _d95, _d96, _d97, _d98, _d99, na3223_93, na3223_94, na3223_95, na3223_96,
                   na3223_97, na3223_98, na3223_99, na3223_100, _d100, _d101, _d102, _d103, _d104, _d105, _d106, _d107, _d108, _d109,
                   _d110, _d111, na3223_113, na3223_114, na3223_115, na3223_116, na3223_117, na3223_118, na3223_119, na3223_120}),
                    .DOBX({_d112, _d113, _d114, _d115, _d116, _d117, _d118, _d119, _d120, _d121, _d122, _d123, _d124, _d125, _d126,
                   _d127, _d128, _d129, _d130, _d131, _d132, _d133, _d134, _d135, _d136, _d137, _d138, _d139, _d140, _d141, _d142, _d143,
                   _d144, _d145, _d146, _d147, _d148, _d149, _d150, _d151}),
                    .ECC1B_ERRA({_d152, _d153, _d154, _d155}),
                    .ECC1B_ERRB({_d156, _d157, _d158, _d159}),
                    .ECC2B_ERRA({_d160, _d161, _d162, _d163}),
                    .ECC2B_ERRB({_d164, _d165, _d166, _d167}),
                    .FORW_CAS_WRAO(_d168), .FORW_CAS_WRBO(_d169), .FORW_CAS_BMAO(_d170), .FORW_CAS_BMBO(_d171), .FORW_CAS_RDAO(_d172),
                    .FORW_CAS_RDBO(_d173), .FORW_UADDRAO({_d174, _d175, _d176, _d177, _d178, _d179, _d180, _d181, _d182, _d183, _d184,
                   _d185, _d186, _d187, _d188, _d189}),
                    .FORW_LADDRAO({_d190, _d191, _d192, _d193, _d194, _d195, _d196, _d197, _d198, _d199, _d200, _d201, _d202, _d203,
                   _d204, _d205}),
                    .FORW_UADDRBO({_d206, _d207, _d208, _d209, _d210, _d211, _d212, _d213, _d214, _d215, _d216, _d217, _d218, _d219,
                   _d220, _d221}),
                    .FORW_LADDRBO({_d222, _d223, _d224, _d225, _d226, _d227, _d228, _d229, _d230, _d231, _d232, _d233, _d234, _d235,
                   _d236, _d237}),
                    .FORW_UA0CLKO(_d238), .FORW_UA0ENO(_d239), .FORW_UA0WEO(_d240), .FORW_LA0CLKO(_d241), .FORW_LA0ENO(_d242), .FORW_LA0WEO(_d243),
                    .FORW_UA1CLKO(_d244), .FORW_UA1ENO(_d245), .FORW_UA1WEO(_d246), .FORW_LA1CLKO(_d247), .FORW_LA1ENO(_d248), .FORW_LA1WEO(_d249),
                    .FORW_UB0CLKO(_d250), .FORW_UB0ENO(_d251), .FORW_UB0WEO(_d252), .FORW_LB0CLKO(_d253), .FORW_LB0ENO(_d254), .FORW_LB0WEO(_d255),
                    .FORW_UB1CLKO(_d256), .FORW_UB1ENO(_d257), .FORW_UB1WEO(_d258), .FORW_LB1CLKO(_d259), .FORW_LB1ENO(_d260), .FORW_LB1WEO(_d261),
                    .CLOCKA({_d262, _d263, _d264, _d265}),
                    .CLOCKB({_d266, _d267, _d268, _d269}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, na3224_10, 1'b1, na3227_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na3232_10, na3233_9, na3236_10, na3237_9, na3238_10, na3239_9, na3240_10, na3242_9, na3244_10, na3245_9,
                   na3250_10, na3251_9, na3253_10, na3257_9, na3261_10, na3264_9}),
                    .ADDRA1({na3265_10, na3266_9, na3269_10, na3271_9, na3273_10, na3277_9, na3280_10, na3284_9, na3286_10, na3289_9,
                   na3291_10, na3293_9, na3294_10, na3295_9, na3297_10, na3299_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({na3300_10, na3304_9, na3306_10, na3308_9, na3309_10, na3311_9, na3314_10, na3315_9, na3318_10, na3319_9,
                   na3320_10, na3321_9, na3323_10, na3325_9, na3326_10, na3330_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({na3332_10, na3333_9, na3337_10, na3339_9, na3340_10, na3344_9, na3345_10, na3347_9, na3349_10, na3350_9,
                   na3351_10, na3352_9, na3353_10, na3354_9, na3355_10, na3356_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na3357_10, na3358_9, na3359_10, na3360_9, na3361_10, na3362_9, na3363_10, na3364_9, na3365_10, na3366_9, 1'b1,
                   1'b1, na3367_10, na3368_9, na3369_10, na3370_9, na3371_10, na3372_9, na3373_10, na3374_9, na3375_10, na3376_9, na3377_10,
                   na3378_9, na3379_10, na3380_9, na3381_10, na3382_9, na3383_10, na3384_9, 1'b1, 1'b1, na3385_10, na3386_9, na3387_10,
                   na3388_9, na3389_10, na3390_9, na3391_10, na3392_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({na3393_10, na3394_9, na3395_10, na3396_9, na3397_10, na3398_9, na3399_10, na3400_9, na3401_10, na3402_9, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na3403_10, na3404_9, na3405_10, na3406_9, na3407_10, na3408_9,
                   na3409_10, na3410_9, na3411_10, na3412_9, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na1739_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
// C_///AND/      x27y41     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3224_4 ( .OUT(na3224_2), .IN1(1'b1), .IN2(na1091_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3224_6 ( .RAM_O2(na3224_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3224_2), .COMP_OUT(1'b0) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_0A_04_00_00_81_03_13_23_00_00_23_00_13_23_00_00_23_00_00),
             .INIT_00(320'h30000014b7000000000000cc50141300000000000000001417000000000000000000130000000000),
             .INIT_01(320'h00015014130000000000000050088300000000000005520023000000000002c70008930000000000),
             .INIT_02(320'h00000088b7000000000000055240230000000000040023889300000000003f802268e30000000000),
             .INIT_03(320'h3f05f3c06f00000000003f802278e300000000003fcf22089300000000001c402208930000000000),
             .INIT_04(320'h080731e46100000000001cc200c83000000000000c0300c0200000000000194721bc430000000000),
             .INIT_05(320'h0000000000000000000000000000000000000000000000286f00000000001b06c194680000000000),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a3225 ( .DOA({_d270, _d271, _d272, _d273, _d274, _d275, _d276, _d277, _d278, _d279, _d280, _d281, _d282, _d283, _d284, _d285,
                   _d286, _d287, _d288, _d289, _d290, _d291, _d292, _d293, _d294, _d295, _d296, _d297, _d298, _d299, _d300, _d301, _d302,
                   _d303, _d304, _d305, _d306, _d307, _d308, _d309}),
                    .DOAX({_d310, _d311, _d312, _d313, _d314, _d315, _d316, _d317, _d318, _d319, _d320, _d321, _d322, _d323, _d324,
                   _d325, _d326, _d327, _d328, _d329, _d330, _d331, _d332, _d333, _d334, _d335, _d336, _d337, _d338, _d339, _d340, _d341,
                   _d342, _d343, _d344, _d345, _d346, _d347, _d348, _d349}),
                    .DOB({_d350, _d351, _d352, _d353, _d354, _d355, _d356, _d357, _d358, _d359, _d360, _d361, na3225_93, na3225_94,
                   na3225_95, na3225_96, na3225_97, na3225_98, na3225_99, na3225_100, _d362, _d363, _d364, _d365, _d366, _d367, _d368,
                   _d369, _d370, _d371, _d372, _d373, _d374, _d375, _d376, _d377, _d378, _d379, _d380, _d381}),
                    .DOBX({_d382, _d383, _d384, _d385, _d386, _d387, _d388, _d389, _d390, _d391, _d392, _d393, _d394, _d395, _d396,
                   _d397, _d398, _d399, _d400, _d401, _d402, _d403, _d404, _d405, _d406, _d407, _d408, _d409, _d410, _d411, _d412, _d413,
                   _d414, _d415, _d416, _d417, _d418, _d419, _d420, _d421}),
                    .ECC1B_ERRA({_d422, _d423, _d424, _d425}),
                    .ECC1B_ERRB({_d426, _d427, _d428, _d429}),
                    .ECC2B_ERRA({_d430, _d431, _d432, _d433}),
                    .ECC2B_ERRB({_d434, _d435, _d436, _d437}),
                    .FORW_CAS_WRAO(_d438), .FORW_CAS_WRBO(_d439), .FORW_CAS_BMAO(_d440), .FORW_CAS_BMBO(_d441), .FORW_CAS_RDAO(_d442),
                    .FORW_CAS_RDBO(_d443), .FORW_UADDRAO({_d444, _d445, _d446, _d447, _d448, _d449, _d450, _d451, _d452, _d453, _d454,
                   _d455, _d456, _d457, _d458, _d459}),
                    .FORW_LADDRAO({_d460, _d461, _d462, _d463, _d464, _d465, _d466, _d467, _d468, _d469, _d470, _d471, _d472, _d473,
                   _d474, _d475}),
                    .FORW_UADDRBO({_d476, _d477, _d478, _d479, _d480, _d481, _d482, _d483, _d484, _d485, _d486, _d487, _d488, _d489,
                   _d490, _d491}),
                    .FORW_LADDRBO({_d492, _d493, _d494, _d495, _d496, _d497, _d498, _d499, _d500, _d501, _d502, _d503, _d504, _d505,
                   _d506, _d507}),
                    .FORW_UA0CLKO(_d508), .FORW_UA0ENO(_d509), .FORW_UA0WEO(_d510), .FORW_LA0CLKO(_d511), .FORW_LA0ENO(_d512), .FORW_LA0WEO(_d513),
                    .FORW_UA1CLKO(_d514), .FORW_UA1ENO(_d515), .FORW_UA1WEO(_d516), .FORW_LA1CLKO(_d517), .FORW_LA1ENO(_d518), .FORW_LA1WEO(_d519),
                    .FORW_UB0CLKO(_d520), .FORW_UB0ENO(_d521), .FORW_UB0WEO(_d522), .FORW_LB0CLKO(_d523), .FORW_LB0ENO(_d524), .FORW_LB0WEO(_d525),
                    .FORW_UB1CLKO(_d526), .FORW_UB1ENO(_d527), .FORW_UB1WEO(_d528), .FORW_LB1CLKO(_d529), .FORW_LB1ENO(_d530), .FORW_LB1WEO(_d531),
                    .CLOCKA({_d532, _d533, _d534, _d535}),
                    .CLOCKB({_d536, _d537, _d538, _d539}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, na3446_10, 1'b1, 1'b1}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1({na3449_10, na3450_9, na3454_10, na3455_9, na3456_10, na3460_9, na3468_10, na3469_9, na3473_10, na3474_9,
                   na3475_10, na3476_9, na3477_10, na3478_9, na3479_10, na3480_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({na3481_10, na3482_9, na3483_10, na3484_9, na3485_10, na3486_9, na3487_10, na3488_9, na3489_10, na3490_9,
                   na3491_10, na3492_9, na3493_10, na3494_9, na3495_10, na3496_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na3497_10, na3498_9, na3499_10, na3500_9, na3501_10, na3502_9, na3503_10, na3504_9, na3505_10, na3506_9, 1'b1,
                   1'b1, na3507_10, na3508_9, na3509_10, na3510_9, na3511_10, na3512_9, na3513_10, na3514_9, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({na3515_10, na3516_9, na3517_10, na3518_9, na3519_10, na3520_9, na3521_10, na3522_9, na3523_10, na3524_9, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na1739_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
FPGA_RAM   #(.RAM_CFG (216'h00_05_00_00_00_00_00_00_0F_04_80_00_91_03_13_23_03_13_23_00_13_23_00_13_23_00_00),
             .INIT_00(320'h30000014b730000014b700cc50141300cc5014130000001417000000141700000000130000000013),
             .INIT_01(320'h00015014130001501413000050088300005008830005520023000552002302c700089302c7000893),
             .INIT_02(320'h00000088b700000088b700055240230005524023040023889304002388933f802268e33f802268e3),
             .INIT_03(320'h3f05f3c06f3f05f3c06f3f802278e33f802278e33fcf2208933fcf2208931c402208931c40220893),
             .INIT_04(320'h080731e461080731e4611cc200d0301cc200cc300c0300c0200c0300c020194721bc43194721bc43),
             .INIT_05(320'h0000000000000000000000000000000000000000000000286f000000286f1b06c194681b06c19468),
             .INIT_06(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_07(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_08(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_09(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_0F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_10(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_11(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_12(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_13(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_14(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_15(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_16(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_17(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_18(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_19(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_1F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_20(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_21(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_22(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_23(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_24(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_25(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_26(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_27(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_28(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_29(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_2F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_30(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_31(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_32(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_33(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_34(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_35(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_36(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_37(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_38(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_39(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_3F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_40(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_41(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_42(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_43(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_44(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_45(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_46(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_47(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_48(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_49(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_4F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_50(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_51(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_52(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_53(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_54(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_55(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_56(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_57(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_58(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_59(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_5F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_60(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_61(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_62(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_63(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_64(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_65(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_66(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_67(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_68(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_69(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_6F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_70(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_71(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_72(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_73(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_74(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_75(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_76(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_77(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_78(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_79(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7A(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7B(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7C(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7D(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7E(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000),
             .INIT_7F(320'h00000000000000000000000000000000000000000000000000000000000000000000000000000000)) 
           _a3226 ( .DOA({_d540, _d541, _d542, _d543, _d544, _d545, _d546, _d547, _d548, _d549, _d550, _d551, _d552, _d553, _d554, _d555,
                   _d556, _d557, _d558, _d559, _d560, _d561, _d562, _d563, _d564, _d565, _d566, _d567, _d568, _d569, _d570, _d571, _d572,
                   _d573, _d574, _d575, _d576, _d577, _d578, _d579}),
                    .DOAX({_d580, _d581, _d582, _d583, _d584, _d585, _d586, _d587, _d588, _d589, _d590, _d591, _d592, _d593, _d594,
                   _d595, _d596, _d597, _d598, _d599, _d600, _d601, _d602, _d603, _d604, _d605, _d606, _d607, _d608, _d609, _d610, _d611,
                   _d612, _d613, _d614, _d615, _d616, _d617, _d618, _d619}),
                    .DOB({_d620, _d621, _d622, _d623, _d624, _d625, _d626, _d627, _d628, _d629, _d630, _d631, na3226_93, na3226_94,
                   na3226_95, na3226_96, na3226_97, na3226_98, na3226_99, na3226_100, _d632, _d633, _d634, _d635, _d636, _d637, _d638,
                   _d639, _d640, _d641, _d642, _d643, na3226_113, na3226_114, na3226_115, na3226_116, na3226_117, na3226_118, na3226_119,
                   na3226_120}),
                    .DOBX({_d644, _d645, _d646, _d647, _d648, _d649, _d650, _d651, _d652, _d653, _d654, _d655, _d656, _d657, _d658,
                   _d659, _d660, _d661, _d662, _d663, _d664, _d665, _d666, _d667, _d668, _d669, _d670, _d671, _d672, _d673, _d674, _d675,
                   _d676, _d677, _d678, _d679, _d680, _d681, _d682, _d683}),
                    .ECC1B_ERRA({_d684, _d685, _d686, _d687}),
                    .ECC1B_ERRB({_d688, _d689, _d690, _d691}),
                    .ECC2B_ERRA({_d692, _d693, _d694, _d695}),
                    .ECC2B_ERRB({_d696, _d697, _d698, _d699}),
                    .FORW_CAS_WRAO(_d700), .FORW_CAS_WRBO(_d701), .FORW_CAS_BMAO(_d702), .FORW_CAS_BMBO(_d703), .FORW_CAS_RDAO(_d704),
                    .FORW_CAS_RDBO(_d705), .FORW_UADDRAO({_d706, _d707, _d708, _d709, _d710, _d711, _d712, _d713, _d714, _d715, _d716,
                   _d717, _d718, _d719, _d720, _d721}),
                    .FORW_LADDRAO({_d722, _d723, _d724, _d725, _d726, _d727, _d728, _d729, _d730, _d731, _d732, _d733, _d734, _d735,
                   _d736, _d737}),
                    .FORW_UADDRBO({_d738, _d739, _d740, _d741, _d742, _d743, _d744, _d745, _d746, _d747, _d748, _d749, _d750, _d751,
                   _d752, _d753}),
                    .FORW_LADDRBO({_d754, _d755, _d756, _d757, _d758, _d759, _d760, _d761, _d762, _d763, _d764, _d765, _d766, _d767,
                   _d768, _d769}),
                    .FORW_UA0CLKO(_d770), .FORW_UA0ENO(_d771), .FORW_UA0WEO(_d772), .FORW_LA0CLKO(_d773), .FORW_LA0ENO(_d774), .FORW_LA0WEO(_d775),
                    .FORW_UA1CLKO(_d776), .FORW_UA1ENO(_d777), .FORW_UA1WEO(_d778), .FORW_LA1CLKO(_d779), .FORW_LA1ENO(_d780), .FORW_LA1WEO(_d781),
                    .FORW_UB0CLKO(_d782), .FORW_UB0ENO(_d783), .FORW_UB0WEO(_d784), .FORW_LB0CLKO(_d785), .FORW_LB0ENO(_d786), .FORW_LB0WEO(_d787),
                    .FORW_UB1CLKO(_d788), .FORW_UB1ENO(_d789), .FORW_UB1WEO(_d790), .FORW_LB1CLKO(_d791), .FORW_LB1ENO(_d792), .FORW_LB1WEO(_d793),
                    .CLOCKA({_d794, _d795, _d796, _d797}),
                    .CLOCKB({_d798, _d799, _d800, _d801}),
                    .CLKA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .CLKB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENA({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ENB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .GLWEA({1'b1, na3533_10, 1'b1, na3534_10}),
                    .GLWEB({1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA0({na3535_10, na3536_9, na3537_10, na3538_9, na3540_10, na3541_9, na3544_10, na3545_9, na3547_10, na3548_9,
                   na3550_10, na3551_9, na3553_10, na3554_9, na3563_10, na3566_9}),
                    .ADDRA1({na3567_10, na3568_9, na3569_10, na3572_9, na3573_10, na3574_9, na3577_10, na3579_9, na3581_10, na3583_9,
                   na3584_10, na3586_9, na3587_10, na3591_9, na3592_10, na3593_9}),
                    .ADDRA0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRA1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB0({na3594_10, na3595_9, na3596_10, na3597_9, na3598_10, na3599_9, na3600_10, na3601_9, na3602_10, na3603_9,
                   na3604_10, na3605_9, na3606_10, na3607_9, na3608_10, na3609_9}),
                    .ADDRB0X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .ADDRB1({na3610_10, na3611_9, na3612_10, na3613_9, na3614_10, na3615_9, na3616_10, na3617_9, na3618_10, na3619_9,
                   na3620_10, na3621_9, na3622_10, na3623_9, na3624_10, na3625_9}),
                    .ADDRB1X({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRA({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .C_ADDRB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .DIA({na3626_10, na3627_9, na3628_10, na3629_9, na3630_10, na3631_9, na3632_10, na3633_9, na3634_10, na3635_9, 1'b1,
                   1'b1, na3636_10, na3637_9, na3638_10, na3639_9, na3640_10, na3641_9, na3642_10, na3643_9, na3644_10, na3645_9, na3646_10,
                   na3647_9, na3648_10, na3649_9, na3650_10, na3651_9, na3652_10, na3653_9, 1'b1, 1'b1, na3654_10, na3655_9, na3656_10,
                   na3658_9, na3659_10, na3662_9, na3663_10, na3665_9}),
                    .DIB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .WEA({na3666_10, na3668_9, na3669_10, na3671_9, na3672_10, na3681_9, na3684_10, na3685_9, na3686_10, na3687_9, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, na3690_10, na3691_9, na3692_10, na3696_9, na3699_10, na3702_9,
                   na3704_10, na3705_9, na3709_10, na3710_9, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .WEB({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1}),
                    .CLOCK1(na1739_1), .CLOCK2(1'b1), .CLOCK3(1'b1), .CLOCK4(1'b1), .FORW_CAS_WRAI(1'b1), .FORW_CAS_WRBI(1'b1), .FORW_CAS_BMAI(1'b1),
                    .FORW_CAS_BMBI(1'b1), .FORW_CAS_RDAI(1'b1), .FORW_CAS_RDBI(1'b1), .FORW_LADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1,
                   1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRAI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_UADDRBI({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
                    .FORW_LA0CLKI(1'b1), .FORW_LA0ENI(1'b1), .FORW_LA0WEI(1'b1), .FORW_UA0CLKI(1'b1), .FORW_UA0ENI(1'b1), .FORW_UA0WEI(1'b1),
                    .FORW_LA1CLKI(1'b1), .FORW_LA1ENI(1'b1), .FORW_LA1WEI(1'b1), .FORW_UA1CLKI(1'b1), .FORW_UA1ENI(1'b1), .FORW_UA1WEI(1'b1),
                    .FORW_LB0CLKI(1'b1), .FORW_LB0ENI(1'b1), .FORW_LB0WEI(1'b1), .FORW_UB0CLKI(1'b1), .FORW_UB0ENI(1'b1), .FORW_UB0WEI(1'b1),
                    .FORW_LB1CLKI(1'b1), .FORW_LB1ENI(1'b1), .FORW_LB1WEI(1'b1), .FORW_UB1CLKI(1'b1), .FORW_UB1ENI(1'b1), .FORW_UB1WEI(1'b1) );
// C_///AND/      x27y33     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3227_4 ( .OUT(na3227_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1233_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3227_6 ( .RAM_O2(na3227_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3227_2), .COMP_OUT(1'b0) );
// C_AND////      x53y63     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3228_1 ( .OUT(na3228_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na709_1), .IN6(1'b1), .IN7(~na2278_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a3229 ( .PCLK0(na3229_1), .PCLK1(na3229_2), .PCLK2(_d802), .PCLK3(_d803), .CLK0(na3219_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0),
                    .SER_CLK(1'b0), .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_///AND/      x52y88     80'h00_0060_00_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3230_4 ( .OUT(na3230_2), .IN1(~na2769_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1050_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x1y128     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3231_5 ( .OUT(na3231_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3222_2), .CP_O(1'b0) );
// C_///AND/      x28y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3232_4 ( .OUT(na3232_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3232_6 ( .RAM_O2(na3232_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3232_2), .COMP_OUT(1'b0) );
// C_AND////      x28y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3233_1 ( .OUT(na3233_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3233_6 ( .RAM_O1(na3233_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3233_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x46y44     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3234_2 ( .OUT(na3234_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3234_6 ( .COUTY1(na3234_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3234_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x13y49     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3235_2 ( .OUT(na3235_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3235_6 ( .COUTY1(na3235_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3235_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3236_4 ( .OUT(na3236_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3236_6 ( .RAM_O2(na3236_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3236_2), .COMP_OUT(1'b0) );
// C_AND////      x28y39     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3237_1 ( .OUT(na3237_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na427_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3237_6 ( .RAM_O1(na3237_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3237_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y38     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3238_4 ( .OUT(na3238_2), .IN1(1'b1), .IN2(na1245_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3238_6 ( .RAM_O2(na3238_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3238_2), .COMP_OUT(1'b0) );
// C_AND////      x28y38     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3239_1 ( .OUT(na3239_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1243_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3239_6 ( .RAM_O1(na3239_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3239_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y37     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3240_4 ( .OUT(na3240_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1241_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3240_6 ( .RAM_O2(na3240_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3240_2), .COMP_OUT(1'b0) );
// C_///AND/      x65y72     80'h00_0060_00_0000_0C08_FF1C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3241_4 ( .OUT(na3241_2), .IN1(1'b1), .IN2(na1986_1), .IN3(~na4485_2), .IN4(~na1990_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y37     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3242_1 ( .OUT(na3242_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1239_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3242_6 ( .RAM_O1(na3242_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3242_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x64y74     80'h00_0018_00_0000_0EEE_3770
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3243_1 ( .OUT(na3243_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na107_1), .IN4(~na104_1), .IN5(~na109_1), .IN6(~na428_1), .IN7(1'b0),
                      .IN8(~na108_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y36     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3244_4 ( .OUT(na3244_2), .IN1(1'b1), .IN2(na1237_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3244_6 ( .RAM_O2(na3244_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3244_2), .COMP_OUT(1'b0) );
// C_AND////      x28y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3245_1 ( .OUT(na3245_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3245_6 ( .RAM_O1(na3245_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3245_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x45y77     80'h00_0018_00_0000_0EEE_C75D
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3246_1 ( .OUT(na3246_1), .IN1(~na984_1), .IN2(na285_2), .IN3(~na83_2), .IN4(1'b0), .IN5(~na1060_1), .IN6(~na12_1), .IN7(1'b0),
                      .IN8(na4153_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x56y65     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3247_2 ( .OUT(na3247_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3247_6 ( .COUTY1(na3247_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3247_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x52y68     80'h00_0018_00_0000_0EEE_7C73
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3248_1 ( .OUT(na3248_1), .IN1(1'b0), .IN2(~na4_1), .IN3(~na83_2), .IN4(~na645_1), .IN5(1'b0), .IN6(na285_1), .IN7(~na736_1),
                      .IN8(~na4154_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y76     80'h00_0018_00_0000_0888_A2C2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3249_1 ( .OUT(na3249_1), .IN1(na1290_1), .IN2(~na285_1), .IN3(1'b1), .IN4(na1208_1), .IN5(na145_1), .IN6(~na285_2), .IN7(na8_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y35     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3250_4 ( .OUT(na3250_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1236_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3250_6 ( .RAM_O2(na3250_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3250_2), .COMP_OUT(1'b0) );
// C_AND////      x28y35     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3251_1 ( .OUT(na3251_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1235_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3251_6 ( .RAM_O1(na3251_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3251_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR////      x16y64     80'h00_0018_00_0000_0C66_C900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3252_1 ( .OUT(na3252_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1483_2), .IN6(~na180_1), .IN7(1'b0), .IN8(na178_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y34     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3253_4 ( .OUT(na3253_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3253_6 ( .RAM_O2(na3253_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3253_2), .COMP_OUT(1'b0) );
// C_///AND/      x16y60     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3254_4 ( .OUT(na3254_2), .IN1(~na2479_2), .IN2(1'b1), .IN3(~na2481_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x17y61     80'h00_0018_00_0000_0888_FC3E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3255_1 ( .OUT(na3255_1), .IN1(na216_1), .IN2(na3258_1), .IN3(1'b0), .IN4(~na3256_2), .IN5(1'b0), .IN6(na3258_2), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x16y58     80'h00_0060_00_0000_0C08_FF75
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3256_4 ( .OUT(na3256_2), .IN1(~na181_1), .IN2(1'b0), .IN3(~na2481_1), .IN4(~na214_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3257_1 ( .OUT(na3257_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3257_6 ( .RAM_O1(na3257_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3257_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND///AND/      x19y60     80'h00_0078_00_0000_0C88_CA58
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3258_1 ( .OUT(na3258_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na216_2), .IN6(1'b1), .IN7(1'b1), .IN8(na214_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3258_4 ( .OUT(na3258_2), .IN1(na4528_2), .IN2(na2478_1), .IN3(~na2481_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x17y47     80'h00_0018_00_0000_0EEE_07C7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3259_1 ( .OUT(na3259_1), .IN1(~na212_1), .IN2(~na209_1), .IN3(1'b0), .IN4(na208_1), .IN5(~na210_1), .IN6(~na1476_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x24y56     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3260_2 ( .OUT(na3260_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3260_6 ( .COUTY1(na3260_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3260_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3261_4 ( .OUT(na3261_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3261_6 ( .RAM_O2(na3261_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3261_2), .COMP_OUT(1'b0) );
// C_MX2b////      x17y46     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3262_1 ( .OUT(na3262_1), .IN1(1'b1), .IN2(na122_1), .IN3(1'b0), .IN4(1'b0), .IN5(na2505_2), .IN6(na132_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x14y59     80'h00_0018_00_0000_0EEE_5733
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3263_1 ( .OUT(na3263_1), .IN1(1'b0), .IN2(~na209_1), .IN3(1'b0), .IN4(~na208_1), .IN5(~na210_1), .IN6(~na1353_1), .IN7(~na211_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3264_1 ( .OUT(na3264_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3264_6 ( .RAM_O1(na3264_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3264_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3265_4 ( .OUT(na3265_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3265_6 ( .RAM_O2(na3265_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3265_2), .COMP_OUT(1'b0) );
// C_AND////      x28y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3266_1 ( .OUT(na3266_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3266_6 ( .RAM_O1(na3266_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3266_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x38y61     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3267_2 ( .OUT(na3267_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3267_6 ( .COUTY1(na3267_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3267_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x20y90     80'h00_0078_00_0000_0C66_0990
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3268_1 ( .OUT(na3268_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2819_2), .IN6(~na387_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3268_4 ( .OUT(na3268_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na388_1), .IN4(na2821_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3269_4 ( .OUT(na3269_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3269_6 ( .RAM_O2(na3269_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3269_2), .COMP_OUT(1'b0) );
// C_///AND/      x46y88     80'h00_0060_00_0000_0C08_FF43
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3270_4 ( .OUT(na3270_2), .IN1(1'b1), .IN2(~na4546_2), .IN3(~na2713_2), .IN4(na2707_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y47     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3271_1 ( .OUT(na3271_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na822_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3271_6 ( .RAM_O1(na3271_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3271_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR////      x60y66     80'h00_0018_00_0000_0C66_6500
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3272_1 ( .OUT(na3272_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na253_1), .IN6(1'b0), .IN7(na251_2), .IN8(na1461_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y46     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3273_4 ( .OUT(na3273_2), .IN1(na1103_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3273_6 ( .RAM_O2(na3273_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3273_2), .COMP_OUT(1'b0) );
// C_///AND/      x57y60     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3274_4 ( .OUT(na3274_2), .IN1(~na2229_1), .IN2(~na2228_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x60y64     80'h00_0018_00_0000_0888_FAE3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3275_1 ( .OUT(na3275_1), .IN1(1'b0), .IN2(~na3276_1), .IN3(na297_1), .IN4(na4583_2), .IN5(na3278_2), .IN6(1'b0), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x57y60     80'h00_0018_00_0000_0C88_57FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3276_1 ( .OUT(na3276_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4512_2), .IN6(~na295_2), .IN7(~na254_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y46     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3277_1 ( .OUT(na3277_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1101_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3277_6 ( .RAM_O1(na3277_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3277_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND///AND/      x57y61     80'h00_0078_00_0000_0C88_ACC4
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3278_1 ( .OUT(na3278_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na295_1), .IN7(na297_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3278_4 ( .OUT(na3278_2), .IN1(~na2229_1), .IN2(na2228_2), .IN3(1'b1), .IN4(na4511_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x31y68     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3279_1 ( .OUT(na3279_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na25_2), .IN7(~na4109_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y45     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3280_4 ( .OUT(na3280_2), .IN1(na1099_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3280_6 ( .RAM_O2(na3280_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3280_2), .COMP_OUT(1'b0) );
// C_/C_0_1///      x62y36     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a3281_2 ( .OUT(na3281_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a3281_6 ( .COUTY1(na3281_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3281_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x52y81     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3282_1 ( .OUT(na3282_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1646_4), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x67y70     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3283_1 ( .OUT(na3283_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1662_4), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y45     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3284_1 ( .OUT(na3284_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1097_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3284_6 ( .RAM_O1(na3284_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3284_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x46y90     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3285_1 ( .OUT(na3285_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1671_4), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y44     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3286_4 ( .OUT(na3286_2), .IN1(1'b1), .IN2(na1095_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3286_6 ( .RAM_O2(na3286_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3286_2), .COMP_OUT(1'b0) );
// C_AND////      x21y59     80'h00_0018_00_0000_0C88_54FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3287_1 ( .OUT(na3287_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na4528_2), .IN6(na2474_1), .IN7(~na4523_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x64y49     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3288_1 ( .OUT(na3288_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1699_4), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y44     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3289_1 ( .OUT(na3289_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3289_6 ( .RAM_O1(na3289_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3289_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND///AND/      x49y71     80'h00_0078_00_0000_0C88_ACAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3290_1 ( .OUT(na3290_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na285_2), .IN7(na139_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3290_4 ( .OUT(na3290_2), .IN1(1'b1), .IN2(na285_1), .IN3(na139_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y43     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3291_4 ( .OUT(na3291_2), .IN1(1'b1), .IN2(na1094_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3291_6 ( .RAM_O2(na3291_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3291_2), .COMP_OUT(1'b0) );
// C_AND////      x22y74     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3292_1 ( .OUT(na3292_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na317_2), .IN8(na4142_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y43     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3293_1 ( .OUT(na3293_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1093_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3293_6 ( .RAM_O1(na3293_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3293_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y42     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3294_4 ( .OUT(na3294_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3294_6 ( .RAM_O2(na3294_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3294_2), .COMP_OUT(1'b0) );
// C_AND////      x28y42     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3295_1 ( .OUT(na3295_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3295_6 ( .RAM_O1(na3295_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3295_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x45y57     80'h00_0078_00_0000_0C66_9090
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3296_1 ( .OUT(na3296_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na713_2), .IN8(~na270_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3296_4 ( .OUT(na3296_2), .IN1(1'b0), .IN2(1'b0), .IN3(na713_1), .IN4(~na270_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y41     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3297_4 ( .OUT(na3297_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3297_6 ( .RAM_O2(na3297_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3297_2), .COMP_OUT(1'b0) );
// C_AND////      x61y57     80'h00_0018_00_0000_0C88_25FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3298_1 ( .OUT(na3298_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2229_2), .IN6(1'b1), .IN7(na2223_1), .IN8(~na4504_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y41     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3299_1 ( .OUT(na3299_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3299_6 ( .RAM_O1(na3299_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3299_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3300_4 ( .OUT(na3300_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3300_6 ( .RAM_O2(na3300_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3300_2), .COMP_OUT(1'b0) );
// C_AND////      x57y70     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3301_1 ( .OUT(na3301_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na349_2), .IN6(~na295_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x68y59     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3302_4 ( .OUT(na3302_2), .IN1(~na351_1), .IN2(1'b0), .IN3(1'b0), .IN4(na4503_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x47y55     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a3303_1 ( .OUT(na3303_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1702_4), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3304_1 ( .OUT(na3304_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3304_6 ( .RAM_O1(na3304_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3304_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x66y48     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3305_4 ( .OUT(na3305_2), .IN1(~na2222_1), .IN2(1'b1), .IN3(~na2223_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3306_4 ( .OUT(na3306_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3306_6 ( .RAM_O2(na3306_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3306_2), .COMP_OUT(1'b0) );
// C_///AND/      x35y81     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3307_4 ( .OUT(na3307_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na287_2), .IN4(na1296_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y39     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3308_1 ( .OUT(na3308_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na427_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3308_6 ( .RAM_O1(na3308_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3308_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y38     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3309_4 ( .OUT(na3309_2), .IN1(1'b1), .IN2(na1288_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3309_6 ( .RAM_O2(na3309_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3309_2), .COMP_OUT(1'b0) );
// C_ORAND////      x22y68     80'h00_0018_00_0000_0C88_B5FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3310_1 ( .OUT(na3310_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na408_1), .IN6(1'b0), .IN7(na4073_2), .IN8(~na27_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y38     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3311_1 ( .OUT(na3311_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1286_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3311_6 ( .RAM_O1(na3311_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3311_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x22y67     80'h00_0018_00_0000_0C88_42FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3312_1 ( .OUT(na3312_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na157_1), .IN6(~na690_1), .IN7(~na11_1), .IN8(na16_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x23y66     80'h00_0018_00_0000_0EEE_57C3
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3313_1 ( .OUT(na3313_1), .IN1(1'b0), .IN2(~na978_1), .IN3(1'b0), .IN4(na926_1), .IN5(~na1520_2), .IN6(~na929_1), .IN7(~na928_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y37     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3314_4 ( .OUT(na3314_2), .IN1(1'b1), .IN2(na1284_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3314_6 ( .RAM_O2(na3314_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3314_2), .COMP_OUT(1'b0) );
// C_AND////      x37y37     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3315_1 ( .OUT(na3315_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1282_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3315_6 ( .RAM_O1(na3315_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3315_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x20y68     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3316_1 ( .OUT(na3316_1), .IN1(1'b1), .IN2(na423_1), .IN3(1'b0), .IN4(1'b0), .IN5(na4579_2), .IN6(na640_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x44y87     80'h00_0018_00_0000_0EEE_7730
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3317_1 ( .OUT(na3317_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(~na409_1), .IN5(~na410_1), .IN6(~na1325_1), .IN7(~na1326_1),
                      .IN8(~na429_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y36     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3318_4 ( .OUT(na3318_2), .IN1(1'b1), .IN2(na1280_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3318_6 ( .RAM_O2(na3318_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3318_2), .COMP_OUT(1'b0) );
// C_AND////      x37y36     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3319_1 ( .OUT(na3319_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3319_6 ( .RAM_O1(na3319_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3319_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y35     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3320_4 ( .OUT(na3320_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1279_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3320_6 ( .RAM_O2(na3320_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3320_2), .COMP_OUT(1'b0) );
// C_AND////      x37y35     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3321_1 ( .OUT(na3321_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1278_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3321_6 ( .RAM_O1(na3321_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3321_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR///XOR/      x63y89     80'h00_0078_00_0000_0C66_0909
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3322_1 ( .OUT(na3322_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1199_2), .IN6(~na1307_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3322_4 ( .OUT(na3322_2), .IN1(na1199_1), .IN2(~na1307_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y34     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3323_4 ( .OUT(na3323_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3323_6 ( .RAM_O2(na3323_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3323_2), .COMP_OUT(1'b0) );
// C_AND////      x60y85     80'h00_0018_00_0000_0C88_A1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3324_1 ( .OUT(na3324_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2962_2), .IN6(~na4566_2), .IN7(na2958_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y34     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3325_1 ( .OUT(na3325_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3325_6 ( .RAM_O1(na3325_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3325_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y33     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3326_4 ( .OUT(na3326_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3326_6 ( .RAM_O2(na3326_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3326_2), .COMP_OUT(1'b0) );
// C_AND////      x49y88     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3327_1 ( .OUT(na3327_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na457_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na4207_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x66y88     80'h00_0060_00_0000_0C06_FFA5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3328_4 ( .OUT(na3328_2), .IN1(~na2957_2), .IN2(1'b0), .IN3(na459_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x62y84     80'h00_0060_00_0000_0C08_FF57
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3329_4 ( .OUT(na3329_2), .IN1(~na456_2), .IN2(~na2965_1), .IN3(~na462_1), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y33     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3330_1 ( .OUT(na3330_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3330_6 ( .RAM_O1(na3330_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3330_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x62y82     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3331_1 ( .OUT(na3331_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2957_2), .IN6(1'b1), .IN7(~na2958_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3332_4 ( .OUT(na3332_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3332_6 ( .RAM_O2(na3332_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3332_2), .COMP_OUT(1'b0) );
// C_AND////      x37y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3333_1 ( .OUT(na3333_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3333_6 ( .RAM_O1(na3333_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3333_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x25y71     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3334_1 ( .OUT(na3334_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na137_2), .IN7(~na3161_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y70     80'h00_0018_00_0000_0C88_ACFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3335_1 ( .OUT(na3335_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na508_2), .IN7(na139_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x65y74     80'h00_0018_00_0000_0C88_75FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3336_1 ( .OUT(na3336_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na513_1), .IN6(1'b0), .IN7(~na38_2), .IN8(~na4492_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3337_4 ( .OUT(na3337_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3337_6 ( .RAM_O2(na3337_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3337_2), .COMP_OUT(1'b0) );
// C_///AND/      x71y69     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3338_4 ( .OUT(na3338_2), .IN1(1'b1), .IN2(~na1986_2), .IN3(1'b1), .IN4(~na1985_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y47     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3339_1 ( .OUT(na3339_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na822_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3339_6 ( .RAM_O1(na3339_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3339_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y46     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3340_4 ( .OUT(na3340_2), .IN1(na1146_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3340_6 ( .RAM_O2(na3340_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3340_2), .COMP_OUT(1'b0) );
// C_ORAND////      x63y70     80'h00_0018_00_0000_0C88_BCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3341_1 ( .OUT(na3341_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na1993_2), .IN7(na4487_2), .IN8(~na1990_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x65y69     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3342_4 ( .OUT(na3342_2), .IN1(1'b1), .IN2(~na1989_2), .IN3(1'b1), .IN4(na1990_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x62y67     80'h00_0018_00_0000_0EEE_57C5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3343_1 ( .OUT(na3343_1), .IN1(~na109_1), .IN2(1'b0), .IN3(1'b0), .IN4(na104_1), .IN5(~na105_1), .IN6(~na1432_1), .IN7(~na107_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y46     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3344_1 ( .OUT(na3344_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1144_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3344_6 ( .RAM_O1(na3344_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3344_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y45     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3345_4 ( .OUT(na3345_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1142_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3345_6 ( .RAM_O2(na3345_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3345_2), .COMP_OUT(1'b0) );
// C_MX2b////      x50y57     80'h00_0018_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3346_1 ( .OUT(na3346_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na55_1), .IN5(1'b0), .IN6(na34_1), .IN7(1'b0), .IN8(na4499_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y45     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3347_1 ( .OUT(na3347_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1140_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3347_6 ( .RAM_O1(na3347_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3347_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_XOR////      x68y75     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3348_1 ( .OUT(na3348_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na522_2), .IN6(1'b0), .IN7(1'b0), .IN8(na1446_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x37y44     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3349_4 ( .OUT(na3349_2), .IN1(1'b1), .IN2(na1138_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3349_6 ( .RAM_O2(na3349_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3349_2), .COMP_OUT(1'b0) );
// C_AND////      x37y44     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3350_1 ( .OUT(na3350_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3350_6 ( .RAM_O1(na3350_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3350_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y43     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3351_4 ( .OUT(na3351_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1137_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3351_6 ( .RAM_O2(na3351_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3351_2), .COMP_OUT(1'b0) );
// C_AND////      x37y43     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3352_1 ( .OUT(na3352_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1136_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3352_6 ( .RAM_O1(na3352_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3352_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y42     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3353_4 ( .OUT(na3353_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3353_6 ( .RAM_O2(na3353_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3353_2), .COMP_OUT(1'b0) );
// C_AND////      x37y42     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3354_1 ( .OUT(na3354_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3354_6 ( .RAM_O1(na3354_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3354_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y41     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3355_4 ( .OUT(na3355_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3355_6 ( .RAM_O2(na3355_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3355_2), .COMP_OUT(1'b0) );
// C_AND////      x37y41     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3356_1 ( .OUT(na3356_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3356_6 ( .RAM_O1(na3356_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3356_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3357_4 ( .OUT(na3357_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3357_6 ( .RAM_O2(na3357_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3357_2), .COMP_OUT(1'b0) );
// C_AND////      x30y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3358_1 ( .OUT(na3358_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3358_6 ( .RAM_O1(na3358_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3358_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3359_4 ( .OUT(na3359_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3359_6 ( .RAM_O2(na3359_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3359_2), .COMP_OUT(1'b0) );
// C_AND////      x30y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3360_1 ( .OUT(na3360_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3360_6 ( .RAM_O1(na3360_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3360_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3361_4 ( .OUT(na3361_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3361_6 ( .RAM_O2(na3361_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3361_2), .COMP_OUT(1'b0) );
// C_AND////      x32y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3362_1 ( .OUT(na3362_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3362_6 ( .RAM_O1(na3362_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3362_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3363_4 ( .OUT(na3363_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3363_6 ( .RAM_O2(na3363_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3363_2), .COMP_OUT(1'b0) );
// C_AND////      x32y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3364_1 ( .OUT(na3364_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3364_6 ( .RAM_O1(na3364_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3364_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y46     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3365_4 ( .OUT(na3365_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3365_6 ( .RAM_O2(na3365_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3365_2), .COMP_OUT(1'b0) );
// C_AND////      x32y46     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3366_1 ( .OUT(na3366_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3366_6 ( .RAM_O1(na3366_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3366_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y44     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3367_4 ( .OUT(na3367_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1135_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3367_6 ( .RAM_O2(na3367_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3367_2), .COMP_OUT(1'b0) );
// C_AND////      x32y44     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3368_1 ( .OUT(na3368_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1111_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3368_6 ( .RAM_O1(na3368_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3368_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y43     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3369_4 ( .OUT(na3369_2), .IN1(1'b1), .IN2(na1110_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3369_6 ( .RAM_O2(na3369_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3369_2), .COMP_OUT(1'b0) );
// C_AND////      x32y43     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3370_1 ( .OUT(na3370_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1109_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3370_6 ( .RAM_O1(na3370_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3370_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y42     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3371_4 ( .OUT(na3371_2), .IN1(na1108_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3371_6 ( .RAM_O2(na3371_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3371_2), .COMP_OUT(1'b0) );
// C_AND////      x32y42     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3372_1 ( .OUT(na3372_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na1107_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3372_6 ( .RAM_O1(na3372_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3372_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y41     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3373_4 ( .OUT(na3373_2), .IN1(na1106_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3373_6 ( .RAM_O2(na3373_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3373_2), .COMP_OUT(1'b0) );
// C_AND////      x32y41     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3374_1 ( .OUT(na3374_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1105_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3374_6 ( .RAM_O1(na3374_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3374_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3375_4 ( .OUT(na3375_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3375_6 ( .RAM_O2(na3375_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3375_2), .COMP_OUT(1'b0) );
// C_AND////      x30y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3376_1 ( .OUT(na3376_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3376_6 ( .RAM_O1(na3376_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3376_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3377_4 ( .OUT(na3377_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3377_6 ( .RAM_O2(na3377_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3377_2), .COMP_OUT(1'b0) );
// C_AND////      x30y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3378_1 ( .OUT(na3378_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3378_6 ( .RAM_O1(na3378_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3378_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3379_4 ( .OUT(na3379_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3379_6 ( .RAM_O2(na3379_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3379_2), .COMP_OUT(1'b0) );
// C_AND////      x32y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3380_1 ( .OUT(na3380_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3380_6 ( .RAM_O1(na3380_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3380_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3381_4 ( .OUT(na3381_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3381_6 ( .RAM_O2(na3381_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3381_2), .COMP_OUT(1'b0) );
// C_AND////      x32y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3382_1 ( .OUT(na3382_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3382_6 ( .RAM_O1(na3382_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3382_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y38     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3383_4 ( .OUT(na3383_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3383_6 ( .RAM_O2(na3383_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3383_2), .COMP_OUT(1'b0) );
// C_AND////      x32y38     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3384_1 ( .OUT(na3384_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3384_6 ( .RAM_O1(na3384_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3384_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y36     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3385_4 ( .OUT(na3385_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1277_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3385_6 ( .RAM_O2(na3385_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3385_2), .COMP_OUT(1'b0) );
// C_AND////      x32y36     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3386_1 ( .OUT(na3386_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1253_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3386_6 ( .RAM_O1(na3386_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3386_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y35     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3387_4 ( .OUT(na3387_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1252_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3387_6 ( .RAM_O2(na3387_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3387_2), .COMP_OUT(1'b0) );
// C_AND////      x32y35     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3388_1 ( .OUT(na3388_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1251_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3388_6 ( .RAM_O1(na3388_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3388_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y34     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3389_4 ( .OUT(na3389_2), .IN1(na1250_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3389_6 ( .RAM_O2(na3389_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3389_2), .COMP_OUT(1'b0) );
// C_AND////      x32y34     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3390_1 ( .OUT(na3390_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1249_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3390_6 ( .RAM_O1(na3390_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3390_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y33     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3391_4 ( .OUT(na3391_2), .IN1(1'b1), .IN2(na1248_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3391_6 ( .RAM_O2(na3391_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3391_2), .COMP_OUT(1'b0) );
// C_AND////      x32y33     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3392_1 ( .OUT(na3392_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na1247_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3392_6 ( .RAM_O1(na3392_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3392_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3393_4 ( .OUT(na3393_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3393_6 ( .RAM_O2(na3393_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3393_2), .COMP_OUT(1'b0) );
// C_AND////      x29y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3394_1 ( .OUT(na3394_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3394_6 ( .RAM_O1(na3394_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3394_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3395_4 ( .OUT(na3395_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3395_6 ( .RAM_O2(na3395_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3395_2), .COMP_OUT(1'b0) );
// C_AND////      x29y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3396_1 ( .OUT(na3396_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3396_6 ( .RAM_O1(na3396_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3396_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y48     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3397_4 ( .OUT(na3397_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3397_6 ( .RAM_O2(na3397_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3397_2), .COMP_OUT(1'b0) );
// C_AND////      x31y48     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3398_1 ( .OUT(na3398_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3398_6 ( .RAM_O1(na3398_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3398_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y47     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3399_4 ( .OUT(na3399_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3399_6 ( .RAM_O2(na3399_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3399_2), .COMP_OUT(1'b0) );
// C_AND////      x31y47     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3400_1 ( .OUT(na3400_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3400_6 ( .RAM_O1(na3400_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3400_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y46     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3401_4 ( .OUT(na3401_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3401_6 ( .RAM_O2(na3401_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3401_2), .COMP_OUT(1'b0) );
// C_AND////      x31y46     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3402_1 ( .OUT(na3402_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3402_6 ( .RAM_O1(na3402_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3402_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3403_4 ( .OUT(na3403_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3403_6 ( .RAM_O2(na3403_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3403_2), .COMP_OUT(1'b0) );
// C_AND////      x29y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3404_1 ( .OUT(na3404_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3404_6 ( .RAM_O1(na3404_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3404_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3405_4 ( .OUT(na3405_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3405_6 ( .RAM_O2(na3405_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3405_2), .COMP_OUT(1'b0) );
// C_AND////      x29y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3406_1 ( .OUT(na3406_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3406_6 ( .RAM_O1(na3406_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3406_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y40     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3407_4 ( .OUT(na3407_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3407_6 ( .RAM_O2(na3407_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3407_2), .COMP_OUT(1'b0) );
// C_AND////      x31y40     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3408_1 ( .OUT(na3408_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3408_6 ( .RAM_O1(na3408_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3408_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y39     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3409_4 ( .OUT(na3409_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3409_6 ( .RAM_O2(na3409_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3409_2), .COMP_OUT(1'b0) );
// C_AND////      x31y39     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3410_1 ( .OUT(na3410_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3410_6 ( .RAM_O1(na3410_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3410_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y38     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3411_4 ( .OUT(na3411_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3411_6 ( .RAM_O2(na3411_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3411_2), .COMP_OUT(1'b0) );
// C_AND////      x31y38     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3412_1 ( .OUT(na3412_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3412_6 ( .RAM_O1(na3412_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3412_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_////RAM_I2      x34y44     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3413_5 ( .OUT(na3413_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_93), .CP_O(1'b0) );
// C_/RAM_I1///      x34y44     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3414_2 ( .OUT(na3414_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_94), .CP_O(1'b0) );
// C_AND////      x70y76     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3415_1 ( .OUT(na3415_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na360_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1985_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x34y43     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3416_5 ( .OUT(na3416_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_95), .CP_O(1'b0) );
// C_/RAM_I1///      x34y43     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3417_2 ( .OUT(na3417_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_96), .CP_O(1'b0) );
// C_AND////      x49y54     80'h00_0018_00_0000_0C88_1FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3418_1 ( .OUT(na3418_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na529_2), .IN8(~na526_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x48y57     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3419_1 ( .OUT(na3419_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na55_1), .IN5(~na48_1), .IN6(1'b0), .IN7(~na2013_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x34y42     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3420_5 ( .OUT(na3420_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_97), .CP_O(1'b0) );
// C_/RAM_I1///      x34y42     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3421_2 ( .OUT(na3421_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_98), .CP_O(1'b0) );
// C_MX2b////      x50y59     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3422_1 ( .OUT(na3422_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na55_1), .IN5(1'b0), .IN6(~na49_1), .IN7(1'b0), .IN8(~na4497_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x34y41     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3423_5 ( .OUT(na3423_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_99), .CP_O(1'b0) );
// C_/RAM_I1///      x34y41     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3424_2 ( .OUT(na3424_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_100), .CP_O(1'b0) );
// C_MX2b////      x56y59     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3425_1 ( .OUT(na3425_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na55_1), .IN5(~na1339_1), .IN6(1'b0), .IN7(~na4498_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x34y36     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3426_5 ( .OUT(na3426_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_113), .CP_O(1'b0) );
// C_/RAM_I1///      x34y36     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3427_2 ( .OUT(na3427_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_114), .CP_O(1'b0) );
// C_MX2b////      x46y59     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3428_1 ( .OUT(na3428_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na55_1), .IN5(1'b0), .IN6(~na44_1), .IN7(1'b0), .IN8(~na2015_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x34y35     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3429_5 ( .OUT(na3429_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_115), .CP_O(1'b0) );
// C_/RAM_I1///      x34y35     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3430_2 ( .OUT(na3430_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_116), .CP_O(1'b0) );
// C_MX2b////      x42y53     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3431_1 ( .OUT(na3431_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na55_1), .IN5(~na45_1), .IN6(1'b0), .IN7(~na2017_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x65y55     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3432_1 ( .OUT(na3432_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2125_1), .IN7(~na529_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y51     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3433_4 ( .OUT(na3433_2), .IN1(1'b1), .IN2(na2125_2), .IN3(~na529_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y50     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3434_4 ( .OUT(na3434_2), .IN1(1'b1), .IN2(na2127_1), .IN3(~na529_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y53     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3435_4 ( .OUT(na3435_2), .IN1(1'b1), .IN2(na2127_2), .IN3(~na529_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x62y58     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3436_1 ( .OUT(na3436_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2129_1), .IN8(~na4224_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x61y60     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3437_1 ( .OUT(na3437_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2129_2), .IN8(~na4224_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x62y61     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3438_1 ( .OUT(na3438_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na529_2), .IN8(na597_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_////RAM_I2      x34y34     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3439_5 ( .OUT(na3439_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_117), .CP_O(1'b0) );
// C_ORAND////      x71y72     80'h00_0018_00_0000_0888_7C5C
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3440_1 ( .OUT(na3440_1), .IN1(1'b0), .IN2(na3453_1), .IN3(~na598_1), .IN4(1'b0), .IN5(1'b0), .IN6(na3453_2), .IN7(~na598_2),
                      .IN8(~na3457_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x63y65     80'h00_0060_00_0000_0C06_FF56
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3441_4 ( .OUT(na3441_2), .IN1(na535_1), .IN2(na599_2), .IN3(~na1447_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/RAM_I1///      x34y34     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3442_2 ( .OUT(na3442_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_118), .CP_O(1'b0) );
// C_////RAM_I2      x34y33     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3443_5 ( .OUT(na3443_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_119), .CP_O(1'b0) );
// C_/RAM_I1///      x34y33     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3444_2 ( .OUT(na3444_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3223_120), .CP_O(1'b0) );
// C_///XOR/      x65y78     80'h00_0060_00_0000_0C06_FF65
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3445_4 ( .OUT(na3445_2), .IN1(~na607_1), .IN2(1'b0), .IN3(na1439_1), .IN4(na605_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x27y9     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3446_4 ( .OUT(na3446_2), .IN1(na930_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3446_6 ( .RAM_O2(na3446_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3446_2), .COMP_OUT(1'b0) );
// C_///AND/      x65y73     80'h00_0060_00_0000_0C08_FF53
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3447_4 ( .OUT(na3447_2), .IN1(1'b1), .IN2(~na1993_2), .IN3(~na1991_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x63y77     80'h00_0018_00_0000_0888_AFE3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3448_1 ( .OUT(na3448_1), .IN1(1'b0), .IN2(~na3336_1), .IN3(na38_1), .IN4(na4603_2), .IN5(1'b1), .IN6(1'b1), .IN7(na3451_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y16     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3449_4 ( .OUT(na3449_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3449_6 ( .RAM_O2(na3449_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3449_2), .COMP_OUT(1'b0) );
// C_AND////      x28y16     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3450_1 ( .OUT(na3450_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3450_6 ( .RAM_O1(na3450_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3450_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND///AND/      x64y75     80'h00_0078_00_0000_0C88_CAC2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3451_1 ( .OUT(na3451_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na360_1), .IN6(1'b1), .IN7(1'b1), .IN8(na4180_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3451_4 ( .OUT(na3451_2), .IN1(na4489_2), .IN2(~na1993_2), .IN3(1'b1), .IN4(na1990_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x65y66     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3452_4 ( .OUT(na3452_2), .IN1(1'b1), .IN2(~na1986_2), .IN3(1'b1), .IN4(na1581_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x69y72     80'h00_0078_00_0000_0CEE_A7D7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3453_1 ( .OUT(na3453_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na619_1), .IN6(~na1986_2), .IN7(na598_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3453_4 ( .OUT(na3453_2), .IN1(~na522_2), .IN2(~na1986_1), .IN3(~na511_2), .IN4(na4486_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y15     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3454_4 ( .OUT(na3454_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3454_6 ( .RAM_O2(na3454_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3454_2), .COMP_OUT(1'b0) );
// C_AND////      x28y15     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3455_1 ( .OUT(na3455_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na198_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3455_6 ( .RAM_O1(na3455_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3455_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y14     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3456_4 ( .OUT(na3456_2), .IN1(1'b1), .IN2(1'b1), .IN3(na942_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3456_6 ( .RAM_O2(na3456_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3456_2), .COMP_OUT(1'b0) );
// C_MX2b////      x68y72     80'h00_0018_00_0040_0AA0_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3457_1 ( .OUT(na3457_1), .IN1(1'b1), .IN2(1'b1), .IN3(na618_1), .IN4(1'b1), .IN5(1'b0), .IN6(na1441_2), .IN7(1'b0), .IN8(na2011_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y57     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3458_4 ( .OUT(na3458_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na529_2), .IN4(na597_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x45y55     80'h00_0018_00_0000_0EEE_50D7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3459_1 ( .OUT(na3459_1), .IN1(~na1387_1), .IN2(~na1383_2), .IN3(~na1454_2), .IN4(na282_1), .IN5(1'b0), .IN6(1'b0), .IN7(~na283_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y14     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3460_1 ( .OUT(na3460_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na940_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3460_6 ( .RAM_O1(na3460_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3460_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x53y56     80'h00_0018_00_0000_0CEE_E000
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3461_1 ( .OUT(na3461_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na276_1), .IN8(na3462_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x52y58     80'h00_0018_00_0000_0888_25C1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3462_1 ( .OUT(na3462_1), .IN1(~na2229_1), .IN2(~na2228_2), .IN3(1'b1), .IN4(na338_2), .IN5(~na2229_2), .IN6(1'b1), .IN7(na332_1),
                      .IN8(~na4432_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x44y51     80'h00_0018_00_0040_0A50_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3463_1 ( .OUT(na3463_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na276_1), .IN4(1'b1), .IN5(na36_1), .IN6(1'b0), .IN7(na4518_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x23y70     80'h00_0018_00_0000_0CEE_3300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3464_1 ( .OUT(na3464_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na137_2), .IN7(1'b0), .IN8(~na3173_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y71     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3465_1 ( .OUT(na3465_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na139_1), .IN8(na645_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x29y69     80'h00_0060_00_0000_0C0E_FF33
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3466_4 ( .OUT(na3466_2), .IN1(1'b0), .IN2(~na137_2), .IN3(1'b0), .IN4(~na3174_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x39y70     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3467_4 ( .OUT(na3467_2), .IN1(1'b1), .IN2(na690_1), .IN3(na139_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y13     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3468_4 ( .OUT(na3468_2), .IN1(1'b1), .IN2(na938_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3468_6 ( .RAM_O2(na3468_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3468_2), .COMP_OUT(1'b0) );
// C_AND////      x28y13     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3469_1 ( .OUT(na3469_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na936_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3469_6 ( .RAM_O1(na3469_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3469_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x62y59     80'h00_0018_00_0000_0C88_BAFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3470_1 ( .OUT(na3470_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2229_1), .IN6(1'b0), .IN7(na2226_2), .IN8(~na4511_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y56     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3471_4 ( .OUT(na3471_2), .IN1(na2229_2), .IN2(1'b1), .IN3(~na2226_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x54y60     80'h00_0018_00_0000_0C66_AA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3472_1 ( .OUT(na3472_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na707_1), .IN6(1'b0), .IN7(na1468_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y12     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3473_4 ( .OUT(na3473_2), .IN1(1'b1), .IN2(1'b1), .IN3(na934_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3473_6 ( .RAM_O2(na3473_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3473_2), .COMP_OUT(1'b0) );
// C_AND////      x28y12     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3474_1 ( .OUT(na3474_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3474_6 ( .RAM_O1(na3474_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3474_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y11     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3475_4 ( .OUT(na3475_2), .IN1(1'b1), .IN2(na933_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3475_6 ( .RAM_O2(na3475_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3475_2), .COMP_OUT(1'b0) );
// C_AND////      x28y11     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3476_1 ( .OUT(na3476_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na932_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3476_6 ( .RAM_O1(na3476_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3476_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y10     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3477_4 ( .OUT(na3477_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3477_6 ( .RAM_O2(na3477_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3477_2), .COMP_OUT(1'b0) );
// C_AND////      x28y10     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3478_1 ( .OUT(na3478_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3478_6 ( .RAM_O1(na3478_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3478_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y9     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3479_4 ( .OUT(na3479_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3479_6 ( .RAM_O2(na3479_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3479_2), .COMP_OUT(1'b0) );
// C_AND////      x28y9     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3480_1 ( .OUT(na3480_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3480_6 ( .RAM_O1(na3480_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3480_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y16     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3481_4 ( .OUT(na3481_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3481_6 ( .RAM_O2(na3481_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3481_2), .COMP_OUT(1'b0) );
// C_AND////      x37y16     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3482_1 ( .OUT(na3482_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3482_6 ( .RAM_O1(na3482_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3482_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y15     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3483_4 ( .OUT(na3483_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3483_6 ( .RAM_O2(na3483_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3483_2), .COMP_OUT(1'b0) );
// C_AND////      x37y15     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3484_1 ( .OUT(na3484_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na198_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3484_6 ( .RAM_O1(na3484_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3484_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y14     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3485_4 ( .OUT(na3485_2), .IN1(na976_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3485_6 ( .RAM_O2(na3485_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3485_2), .COMP_OUT(1'b0) );
// C_AND////      x37y14     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3486_1 ( .OUT(na3486_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na974_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3486_6 ( .RAM_O1(na3486_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3486_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y13     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3487_4 ( .OUT(na3487_2), .IN1(1'b1), .IN2(1'b1), .IN3(na972_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3487_6 ( .RAM_O2(na3487_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3487_2), .COMP_OUT(1'b0) );
// C_AND////      x37y13     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3488_1 ( .OUT(na3488_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na970_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3488_6 ( .RAM_O1(na3488_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3488_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y12     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3489_4 ( .OUT(na3489_2), .IN1(1'b1), .IN2(na968_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3489_6 ( .RAM_O2(na3489_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3489_2), .COMP_OUT(1'b0) );
// C_AND////      x37y12     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3490_1 ( .OUT(na3490_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3490_6 ( .RAM_O1(na3490_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3490_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y11     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3491_4 ( .OUT(na3491_2), .IN1(1'b1), .IN2(na967_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3491_6 ( .RAM_O2(na3491_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3491_2), .COMP_OUT(1'b0) );
// C_AND////      x37y11     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3492_1 ( .OUT(na3492_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na966_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3492_6 ( .RAM_O1(na3492_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3492_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y10     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3493_4 ( .OUT(na3493_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3493_6 ( .RAM_O2(na3493_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3493_2), .COMP_OUT(1'b0) );
// C_AND////      x37y10     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3494_1 ( .OUT(na3494_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3494_6 ( .RAM_O1(na3494_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3494_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y9     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3495_4 ( .OUT(na3495_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3495_6 ( .RAM_O2(na3495_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3495_2), .COMP_OUT(1'b0) );
// C_AND////      x37y9     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3496_1 ( .OUT(na3496_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3496_6 ( .RAM_O1(na3496_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3496_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y16     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3497_4 ( .OUT(na3497_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3497_6 ( .RAM_O2(na3497_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3497_2), .COMP_OUT(1'b0) );
// C_AND////      x30y16     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3498_1 ( .OUT(na3498_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3498_6 ( .RAM_O1(na3498_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3498_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y15     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3499_4 ( .OUT(na3499_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3499_6 ( .RAM_O2(na3499_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3499_2), .COMP_OUT(1'b0) );
// C_AND////      x30y15     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3500_1 ( .OUT(na3500_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3500_6 ( .RAM_O1(na3500_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3500_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y16     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3501_4 ( .OUT(na3501_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3501_6 ( .RAM_O2(na3501_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3501_2), .COMP_OUT(1'b0) );
// C_AND////      x32y16     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3502_1 ( .OUT(na3502_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3502_6 ( .RAM_O1(na3502_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3502_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y15     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3503_4 ( .OUT(na3503_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3503_6 ( .RAM_O2(na3503_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3503_2), .COMP_OUT(1'b0) );
// C_AND////      x32y15     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3504_1 ( .OUT(na3504_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3504_6 ( .RAM_O1(na3504_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3504_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y14     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3505_4 ( .OUT(na3505_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3505_6 ( .RAM_O2(na3505_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3505_2), .COMP_OUT(1'b0) );
// C_AND////      x32y14     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3506_1 ( .OUT(na3506_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3506_6 ( .RAM_O1(na3506_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3506_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y12     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3507_4 ( .OUT(na3507_2), .IN1(na965_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3507_6 ( .RAM_O2(na3507_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3507_2), .COMP_OUT(1'b0) );
// C_AND////      x32y12     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3508_1 ( .OUT(na3508_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na950_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3508_6 ( .RAM_O1(na3508_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3508_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y11     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3509_4 ( .OUT(na3509_2), .IN1(na949_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3509_6 ( .RAM_O2(na3509_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3509_2), .COMP_OUT(1'b0) );
// C_AND////      x32y11     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3510_1 ( .OUT(na3510_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na948_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3510_6 ( .RAM_O1(na3510_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3510_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y10     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3511_4 ( .OUT(na3511_2), .IN1(1'b1), .IN2(1'b1), .IN3(na947_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3511_6 ( .RAM_O2(na3511_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3511_2), .COMP_OUT(1'b0) );
// C_AND////      x32y10     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3512_1 ( .OUT(na3512_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na946_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3512_6 ( .RAM_O1(na3512_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3512_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y9     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3513_4 ( .OUT(na3513_2), .IN1(na945_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3513_6 ( .RAM_O2(na3513_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3513_2), .COMP_OUT(1'b0) );
// C_AND////      x32y9     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3514_1 ( .OUT(na3514_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na944_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3514_6 ( .RAM_O1(na3514_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3514_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y16     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3515_4 ( .OUT(na3515_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3515_6 ( .RAM_O2(na3515_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3515_2), .COMP_OUT(1'b0) );
// C_AND////      x29y16     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3516_1 ( .OUT(na3516_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3516_6 ( .RAM_O1(na3516_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3516_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y15     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3517_4 ( .OUT(na3517_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3517_6 ( .RAM_O2(na3517_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3517_2), .COMP_OUT(1'b0) );
// C_AND////      x29y15     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3518_1 ( .OUT(na3518_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3518_6 ( .RAM_O1(na3518_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3518_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y16     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3519_4 ( .OUT(na3519_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3519_6 ( .RAM_O2(na3519_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3519_2), .COMP_OUT(1'b0) );
// C_AND////      x31y16     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3520_1 ( .OUT(na3520_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3520_6 ( .RAM_O1(na3520_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3520_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y15     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3521_4 ( .OUT(na3521_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3521_6 ( .RAM_O2(na3521_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3521_2), .COMP_OUT(1'b0) );
// C_AND////      x31y15     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3522_1 ( .OUT(na3522_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3522_6 ( .RAM_O1(na3522_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3522_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y14     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3523_4 ( .OUT(na3523_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3523_6 ( .RAM_O2(na3523_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3523_2), .COMP_OUT(1'b0) );
// C_AND////      x31y14     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3524_1 ( .OUT(na3524_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3524_6 ( .RAM_O1(na3524_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3524_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_////RAM_I2      x34y12     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3525_5 ( .OUT(na3525_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3225_93), .CP_O(1'b0) );
// C_/RAM_I1///      x34y12     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3526_2 ( .OUT(na3526_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3225_94), .CP_O(1'b0) );
// C_////RAM_I2      x34y11     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3527_5 ( .OUT(na3527_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3225_95), .CP_O(1'b0) );
// C_/RAM_I1///      x34y11     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3528_2 ( .OUT(na3528_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3225_96), .CP_O(1'b0) );
// C_////RAM_I2      x34y10     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3529_5 ( .OUT(na3529_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3225_97), .CP_O(1'b0) );
// C_/RAM_I1///      x34y10     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3530_2 ( .OUT(na3530_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3225_98), .CP_O(1'b0) );
// C_////RAM_I2      x34y9     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3531_5 ( .OUT(na3531_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3225_99), .CP_O(1'b0) );
// C_/RAM_I1///      x34y9     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3532_2 ( .OUT(na3532_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3225_100), .CP_O(1'b0) );
// C_///AND/      x27y25     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3533_4 ( .OUT(na3533_2), .IN1(1'b1), .IN2(1'b1), .IN3(na576_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3533_6 ( .RAM_O2(na3533_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3533_2), .COMP_OUT(1'b0) );
// C_///AND/      x27y17     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3534_4 ( .OUT(na3534_2), .IN1(na763_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3534_6 ( .RAM_O2(na3534_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3534_2), .COMP_OUT(1'b0) );
// C_///AND/      x28y24     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3535_4 ( .OUT(na3535_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3535_6 ( .RAM_O2(na3535_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3535_2), .COMP_OUT(1'b0) );
// C_AND////      x28y24     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3536_1 ( .OUT(na3536_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3536_6 ( .RAM_O1(na3536_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3536_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y23     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3537_4 ( .OUT(na3537_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3537_6 ( .RAM_O2(na3537_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3537_2), .COMP_OUT(1'b0) );
// C_AND////      x28y23     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3538_1 ( .OUT(na3538_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na639_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3538_6 ( .RAM_O1(na3538_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3538_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x65y58     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3539_1 ( .OUT(na3539_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2222_1), .IN6(1'b1), .IN7(na297_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y22     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3540_4 ( .OUT(na3540_2), .IN1(1'b1), .IN2(1'b1), .IN3(na775_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3540_6 ( .RAM_O2(na3540_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3540_2), .COMP_OUT(1'b0) );
// C_AND////      x28y22     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3541_1 ( .OUT(na3541_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na773_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3541_6 ( .RAM_O1(na3541_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3541_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x49y47     80'h00_0018_00_0000_0C88_55FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3542_1 ( .OUT(na3542_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na638_2), .IN6(1'b1), .IN7(~na636_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x48y54     80'h00_0018_00_0040_0A55_00A0
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3543_1 ( .OUT(na3543_1), .IN1(1'b0), .IN2(1'b0), .IN3(na276_1), .IN4(1'b1), .IN5(~na2250_1), .IN6(1'b0), .IN7(~na323_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y21     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3544_4 ( .OUT(na3544_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na771_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3544_6 ( .RAM_O2(na3544_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3544_2), .COMP_OUT(1'b0) );
// C_AND////      x28y21     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3545_1 ( .OUT(na3545_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na769_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3545_6 ( .RAM_O1(na3545_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3545_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x48y56     80'h00_0018_00_0040_0AAA_00AF
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3546_1 ( .OUT(na3546_1), .IN1(1'b1), .IN2(1'b1), .IN3(na276_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na4516_2), .IN7(1'b0), .IN8(~na162_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y20     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3547_4 ( .OUT(na3547_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na767_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3547_6 ( .RAM_O2(na3547_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3547_2), .COMP_OUT(1'b0) );
// C_AND////      x28y20     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3548_1 ( .OUT(na3548_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3548_6 ( .RAM_O1(na3548_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3548_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x48y52     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3549_1 ( .OUT(na3549_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na276_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na324_1), .IN7(1'b0), .IN8(~na4517_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y19     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3550_4 ( .OUT(na3550_2), .IN1(1'b1), .IN2(1'b1), .IN3(na766_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3550_6 ( .RAM_O2(na3550_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3550_2), .COMP_OUT(1'b0) );
// C_AND////      x28y19     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3551_1 ( .OUT(na3551_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na765_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3551_6 ( .RAM_O1(na3551_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3551_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x44y52     80'h00_0018_00_0040_0A55_0050
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3552_1 ( .OUT(na3552_1), .IN1(1'b0), .IN2(1'b0), .IN3(~na276_1), .IN4(1'b1), .IN5(~na325_1), .IN6(1'b0), .IN7(~na2252_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y18     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3553_4 ( .OUT(na3553_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3553_6 ( .RAM_O2(na3553_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3553_2), .COMP_OUT(1'b0) );
// C_AND////      x28y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3554_1 ( .OUT(na3554_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3554_6 ( .RAM_O1(na3554_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3554_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x42y52     80'h00_0018_00_0040_0AAA_005F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3555_1 ( .OUT(na3555_1), .IN1(1'b1), .IN2(1'b1), .IN3(~na276_1), .IN4(1'b1), .IN5(1'b0), .IN6(~na315_1), .IN7(1'b0), .IN8(~na2254_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x59y41     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3556_4 ( .OUT(na3556_2), .IN1(~na638_2), .IN2(na2359_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y42     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3557_4 ( .OUT(na3557_2), .IN1(~na638_2), .IN2(na2359_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x57y41     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3558_4 ( .OUT(na3558_2), .IN1(~na638_2), .IN2(1'b1), .IN3(na2361_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x57y44     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3559_1 ( .OUT(na3559_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na638_2), .IN6(1'b1), .IN7(na2361_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x58y41     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3560_1 ( .OUT(na3560_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na638_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2363_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x61y44     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3561_1 ( .OUT(na3561_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na638_2), .IN6(1'b1), .IN7(1'b1), .IN8(na2363_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x51y43     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3562_4 ( .OUT(na3562_2), .IN1(~na638_2), .IN2(1'b1), .IN3(na784_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3563_4 ( .OUT(na3563_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3563_6 ( .RAM_O2(na3563_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3563_2), .COMP_OUT(1'b0) );
// C_ORAND////      x67y57     80'h00_0018_00_0000_0888_A7A5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3564_1 ( .OUT(na3564_1), .IN1(~na785_1), .IN2(1'b0), .IN3(na3571_1), .IN4(1'b0), .IN5(~na785_2), .IN6(~na3575_1), .IN7(na3571_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x61y50     80'h00_0060_00_0000_0C06_FF9C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3565_4 ( .OUT(na3565_2), .IN1(1'b0), .IN2(na786_1), .IN3(~na1469_1), .IN4(na720_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3566_1 ( .OUT(na3566_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3566_6 ( .RAM_O1(na3566_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3566_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y32     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3567_4 ( .OUT(na3567_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3567_6 ( .RAM_O2(na3567_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3567_2), .COMP_OUT(1'b0) );
// C_AND////      x28y32     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3568_1 ( .OUT(na3568_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3568_6 ( .RAM_O1(na3568_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3568_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y31     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3569_4 ( .OUT(na3569_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3569_6 ( .RAM_O2(na3569_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3569_2), .COMP_OUT(1'b0) );
// C_///AND/      x61y47     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3570_4 ( .OUT(na3570_2), .IN1(1'b1), .IN2(na1587_2), .IN3(~na2223_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x68y55     80'h00_0078_00_0000_0CEE_7AD7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3571_1 ( .OUT(na3571_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na785_2), .IN6(1'b0), .IN7(~na797_1), .IN8(~na4504_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3571_4 ( .OUT(na3571_2), .IN1(~na707_1), .IN2(~na352_2), .IN3(~na2223_1), .IN4(na4504_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y31     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3572_1 ( .OUT(na3572_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na530_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3572_6 ( .RAM_O1(na3572_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3572_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y30     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3573_4 ( .OUT(na3573_2), .IN1(na588_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3573_6 ( .RAM_O2(na3573_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3573_2), .COMP_OUT(1'b0) );
// C_AND////      x28y30     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3574_1 ( .OUT(na3574_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na586_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3574_6 ( .RAM_O1(na3574_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3574_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_MX2b////      x61y56     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3575_1 ( .OUT(na3575_1), .IN1(1'b1), .IN2(na796_2), .IN3(1'b0), .IN4(1'b0), .IN5(na1463_1), .IN6(na2248_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x55y53     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3576_4 ( .OUT(na3576_2), .IN1(~na638_2), .IN2(1'b1), .IN3(na784_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y29     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3577_4 ( .OUT(na3577_2), .IN1(1'b1), .IN2(1'b1), .IN3(na584_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3577_6 ( .RAM_O2(na3577_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3577_2), .COMP_OUT(1'b0) );
// C_OR////      x41y85     80'h00_0018_00_0000_0EEE_55C7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3578_1 ( .OUT(na3578_1), .IN1(~na1498_1), .IN2(~na1325_1), .IN3(1'b0), .IN4(na409_1), .IN5(~na430_2), .IN6(1'b0), .IN7(~na1326_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y29     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3579_1 ( .OUT(na3579_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na582_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3579_6 ( .RAM_O1(na3579_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3579_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_OR////      x40y81     80'h00_0018_00_0000_0EEE_7EAC
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3580_1 ( .OUT(na3580_1), .IN1(1'b0), .IN2(na4553_2), .IN3(na2713_1), .IN4(1'b0), .IN5(na2712_2), .IN6(na232_1), .IN7(~na1340_1),
                      .IN8(~na3230_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x28y28     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3581_4 ( .OUT(na3581_2), .IN1(1'b1), .IN2(na580_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3581_6 ( .RAM_O2(na3581_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3581_2), .COMP_OUT(1'b0) );
// C_MX2b////      x30y72     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3582_1 ( .OUT(na3582_1), .IN1(1'b1), .IN2(na219_2), .IN3(1'b0), .IN4(1'b0), .IN5(na4561_2), .IN6(na1312_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y28     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3583_1 ( .OUT(na3583_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3583_6 ( .RAM_O1(na3583_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3583_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y27     80'h08_0060_00_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3584_4 ( .OUT(na3584_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na579_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3584_6 ( .RAM_O2(na3584_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3584_2), .COMP_OUT(1'b0) );
// C_AND////      x27y57     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3585_1 ( .OUT(na3585_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2474_2), .IN7(1'b1), .IN8(~na2473_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y27     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3586_1 ( .OUT(na3586_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na578_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3586_6 ( .RAM_O1(na3586_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3586_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y26     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3587_4 ( .OUT(na3587_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3587_6 ( .RAM_O2(na3587_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3587_2), .COMP_OUT(1'b0) );
// C_ORAND////      x22y57     80'h00_0018_00_0000_0C88_ABFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3588_1 ( .OUT(na3588_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4524_2), .IN6(~na2478_2), .IN7(na2481_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x22y54     80'h00_0018_00_0000_0C88_F2FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3589_1 ( .OUT(na3589_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na4530_2), .IN6(~na2477_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x15y53     80'h00_0018_00_0000_0C66_CA00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3590_1 ( .OUT(na3590_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1490_2), .IN6(1'b0), .IN7(1'b0), .IN8(na884_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x28y26     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3591_1 ( .OUT(na3591_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3591_6 ( .RAM_O1(na3591_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3591_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x28y25     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3592_4 ( .OUT(na3592_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3592_6 ( .RAM_O2(na3592_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3592_2), .COMP_OUT(1'b0) );
// C_AND////      x28y25     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3593_1 ( .OUT(na3593_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3593_6 ( .RAM_O1(na3593_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3593_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y24     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3594_4 ( .OUT(na3594_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3594_6 ( .RAM_O2(na3594_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3594_2), .COMP_OUT(1'b0) );
// C_AND////      x37y24     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3595_1 ( .OUT(na3595_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3595_6 ( .RAM_O1(na3595_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3595_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y23     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3596_4 ( .OUT(na3596_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3596_6 ( .RAM_O2(na3596_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3596_2), .COMP_OUT(1'b0) );
// C_AND////      x37y23     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3597_1 ( .OUT(na3597_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na639_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3597_6 ( .RAM_O1(na3597_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3597_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y22     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3598_4 ( .OUT(na3598_2), .IN1(1'b1), .IN2(1'b1), .IN3(na809_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3598_6 ( .RAM_O2(na3598_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3598_2), .COMP_OUT(1'b0) );
// C_AND////      x37y22     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3599_1 ( .OUT(na3599_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na807_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3599_6 ( .RAM_O1(na3599_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3599_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y21     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3600_4 ( .OUT(na3600_2), .IN1(na805_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3600_6 ( .RAM_O2(na3600_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3600_2), .COMP_OUT(1'b0) );
// C_AND////      x37y21     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3601_1 ( .OUT(na3601_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na803_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3601_6 ( .RAM_O1(na3601_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3601_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y20     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3602_4 ( .OUT(na3602_2), .IN1(na801_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3602_6 ( .RAM_O2(na3602_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3602_2), .COMP_OUT(1'b0) );
// C_AND////      x37y20     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3603_1 ( .OUT(na3603_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3603_6 ( .RAM_O1(na3603_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3603_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y19     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3604_4 ( .OUT(na3604_2), .IN1(1'b1), .IN2(1'b1), .IN3(na800_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3604_6 ( .RAM_O2(na3604_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3604_2), .COMP_OUT(1'b0) );
// C_AND////      x37y19     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3605_1 ( .OUT(na3605_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na799_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3605_6 ( .RAM_O1(na3605_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3605_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y18     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3606_4 ( .OUT(na3606_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3606_6 ( .RAM_O2(na3606_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3606_2), .COMP_OUT(1'b0) );
// C_AND////      x37y18     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3607_1 ( .OUT(na3607_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3607_6 ( .RAM_O1(na3607_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3607_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y17     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3608_4 ( .OUT(na3608_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3608_6 ( .RAM_O2(na3608_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3608_2), .COMP_OUT(1'b0) );
// C_AND////      x37y17     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3609_1 ( .OUT(na3609_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3609_6 ( .RAM_O1(na3609_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3609_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y32     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3610_4 ( .OUT(na3610_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3610_6 ( .RAM_O2(na3610_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3610_2), .COMP_OUT(1'b0) );
// C_AND////      x37y32     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3611_1 ( .OUT(na3611_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3611_6 ( .RAM_O1(na3611_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3611_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y31     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3612_4 ( .OUT(na3612_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3612_6 ( .RAM_O2(na3612_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3612_2), .COMP_OUT(1'b0) );
// C_AND////      x37y31     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3613_1 ( .OUT(na3613_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na530_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3613_6 ( .RAM_O1(na3613_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3613_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y30     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3614_4 ( .OUT(na3614_2), .IN1(1'b1), .IN2(na631_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3614_6 ( .RAM_O2(na3614_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3614_2), .COMP_OUT(1'b0) );
// C_AND////      x37y30     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3615_1 ( .OUT(na3615_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na629_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3615_6 ( .RAM_O1(na3615_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3615_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y29     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3616_4 ( .OUT(na3616_2), .IN1(1'b1), .IN2(1'b1), .IN3(na627_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3616_6 ( .RAM_O2(na3616_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3616_2), .COMP_OUT(1'b0) );
// C_AND////      x37y29     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3617_1 ( .OUT(na3617_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na625_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3617_6 ( .RAM_O1(na3617_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3617_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y28     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3618_4 ( .OUT(na3618_2), .IN1(na623_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3618_6 ( .RAM_O2(na3618_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3618_2), .COMP_OUT(1'b0) );
// C_AND////      x37y28     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3619_1 ( .OUT(na3619_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3619_6 ( .RAM_O1(na3619_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3619_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y27     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3620_4 ( .OUT(na3620_2), .IN1(na622_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3620_6 ( .RAM_O2(na3620_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3620_2), .COMP_OUT(1'b0) );
// C_AND////      x37y27     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3621_1 ( .OUT(na3621_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na621_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3621_6 ( .RAM_O1(na3621_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3621_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y26     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3622_4 ( .OUT(na3622_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3622_6 ( .RAM_O2(na3622_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3622_2), .COMP_OUT(1'b0) );
// C_AND////      x37y26     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3623_1 ( .OUT(na3623_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3623_6 ( .RAM_O1(na3623_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3623_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y25     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3624_4 ( .OUT(na3624_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3624_6 ( .RAM_O2(na3624_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3624_2), .COMP_OUT(1'b0) );
// C_AND////      x37y25     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3625_1 ( .OUT(na3625_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3625_6 ( .RAM_O1(na3625_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3625_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y32     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3626_4 ( .OUT(na3626_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3626_6 ( .RAM_O2(na3626_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3626_2), .COMP_OUT(1'b0) );
// C_AND////      x30y32     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3627_1 ( .OUT(na3627_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3627_6 ( .RAM_O1(na3627_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3627_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y31     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3628_4 ( .OUT(na3628_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3628_6 ( .RAM_O2(na3628_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3628_2), .COMP_OUT(1'b0) );
// C_AND////      x30y31     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3629_1 ( .OUT(na3629_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3629_6 ( .RAM_O1(na3629_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3629_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y32     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3630_4 ( .OUT(na3630_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3630_6 ( .RAM_O2(na3630_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3630_2), .COMP_OUT(1'b0) );
// C_AND////      x32y32     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3631_1 ( .OUT(na3631_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3631_6 ( .RAM_O1(na3631_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3631_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y31     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3632_4 ( .OUT(na3632_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3632_6 ( .RAM_O2(na3632_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3632_2), .COMP_OUT(1'b0) );
// C_AND////      x32y31     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3633_1 ( .OUT(na3633_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3633_6 ( .RAM_O1(na3633_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3633_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y30     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3634_4 ( .OUT(na3634_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3634_6 ( .RAM_O2(na3634_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3634_2), .COMP_OUT(1'b0) );
// C_AND////      x32y30     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3635_1 ( .OUT(na3635_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3635_6 ( .RAM_O1(na3635_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3635_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y28     80'h08_0060_00_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3636_4 ( .OUT(na3636_2), .IN1(1'b1), .IN2(na620_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3636_6 ( .RAM_O2(na3636_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3636_2), .COMP_OUT(1'b0) );
// C_AND////      x32y28     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3637_1 ( .OUT(na3637_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na596_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3637_6 ( .RAM_O1(na3637_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3637_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y27     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3638_4 ( .OUT(na3638_2), .IN1(1'b1), .IN2(1'b1), .IN3(na595_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3638_6 ( .RAM_O2(na3638_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3638_2), .COMP_OUT(1'b0) );
// C_AND////      x32y27     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3639_1 ( .OUT(na3639_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na594_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3639_6 ( .RAM_O1(na3639_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3639_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y26     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3640_4 ( .OUT(na3640_2), .IN1(na593_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3640_6 ( .RAM_O2(na3640_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3640_2), .COMP_OUT(1'b0) );
// C_AND////      x32y26     80'h04_0018_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3641_1 ( .OUT(na3641_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na592_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3641_6 ( .RAM_O1(na3641_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3641_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y25     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3642_4 ( .OUT(na3642_2), .IN1(1'b1), .IN2(1'b1), .IN3(na591_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3642_6 ( .RAM_O2(na3642_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3642_2), .COMP_OUT(1'b0) );
// C_AND////      x32y25     80'h04_0018_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3643_1 ( .OUT(na3643_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na590_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3643_6 ( .RAM_O1(na3643_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3643_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y24     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3644_4 ( .OUT(na3644_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3644_6 ( .RAM_O2(na3644_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3644_2), .COMP_OUT(1'b0) );
// C_AND////      x30y24     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3645_1 ( .OUT(na3645_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3645_6 ( .RAM_O1(na3645_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3645_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x30y23     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3646_4 ( .OUT(na3646_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3646_6 ( .RAM_O2(na3646_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3646_2), .COMP_OUT(1'b0) );
// C_AND////      x30y23     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3647_1 ( .OUT(na3647_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3647_6 ( .RAM_O1(na3647_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3647_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y24     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3648_4 ( .OUT(na3648_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3648_6 ( .RAM_O2(na3648_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3648_2), .COMP_OUT(1'b0) );
// C_AND////      x32y24     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3649_1 ( .OUT(na3649_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3649_6 ( .RAM_O1(na3649_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3649_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y23     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3650_4 ( .OUT(na3650_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3650_6 ( .RAM_O2(na3650_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3650_2), .COMP_OUT(1'b0) );
// C_AND////      x32y23     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3651_1 ( .OUT(na3651_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3651_6 ( .RAM_O1(na3651_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3651_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y22     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3652_4 ( .OUT(na3652_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3652_6 ( .RAM_O2(na3652_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3652_2), .COMP_OUT(1'b0) );
// C_AND////      x32y22     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3653_1 ( .OUT(na3653_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3653_6 ( .RAM_O1(na3653_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3653_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y20     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3654_4 ( .OUT(na3654_2), .IN1(na798_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3654_6 ( .RAM_O2(na3654_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3654_2), .COMP_OUT(1'b0) );
// C_AND////      x32y20     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3655_1 ( .OUT(na3655_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na783_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3655_6 ( .RAM_O1(na3655_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3655_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y19     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3656_4 ( .OUT(na3656_2), .IN1(1'b1), .IN2(1'b1), .IN3(na782_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3656_6 ( .RAM_O2(na3656_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3656_2), .COMP_OUT(1'b0) );
// C_///AND/      x30y62     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3657_4 ( .OUT(na3657_2), .IN1(na216_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2473_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x32y19     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3658_1 ( .OUT(na3658_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na781_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3658_6 ( .RAM_O1(na3658_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3658_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y18     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3659_4 ( .OUT(na3659_2), .IN1(na780_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3659_6 ( .RAM_O2(na3659_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3659_2), .COMP_OUT(1'b0) );
// C_///AND/      x14y47     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3660_4 ( .OUT(na3660_2), .IN1(1'b1), .IN2(~na194_1), .IN3(1'b1), .IN4(~na197_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x19y43     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3661_1 ( .OUT(na3661_1), .IN1(1'b1), .IN2(na122_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2501_1), .IN6(~na126_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x32y18     80'h04_0018_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3662_1 ( .OUT(na3662_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na779_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3662_6 ( .RAM_O1(na3662_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3662_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x32y17     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3663_4 ( .OUT(na3663_2), .IN1(1'b1), .IN2(1'b1), .IN3(na778_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3663_6 ( .RAM_O2(na3663_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3663_2), .COMP_OUT(1'b0) );
// C_MX2b////      x21y43     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3664_1 ( .OUT(na3664_1), .IN1(1'b1), .IN2(~na122_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1367_1), .IN6(~na4539_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x32y17     80'h04_0018_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3665_1 ( .OUT(na3665_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na777_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3665_6 ( .RAM_O1(na3665_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3665_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y32     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3666_4 ( .OUT(na3666_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3666_6 ( .RAM_O2(na3666_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3666_2), .COMP_OUT(1'b0) );
// C_MX2b////      x17y41     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3667_1 ( .OUT(na3667_1), .IN1(1'b1), .IN2(~na122_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1366_1), .IN6(~na2503_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y32     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3668_1 ( .OUT(na3668_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3668_6 ( .RAM_O1(na3668_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3668_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y31     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3669_4 ( .OUT(na3669_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3669_6 ( .RAM_O2(na3669_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3669_2), .COMP_OUT(1'b0) );
// C_MX2b////      x17y43     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3670_1 ( .OUT(na3670_1), .IN1(1'b1), .IN2(na122_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na4540_2), .IN6(~na130_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y31     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3671_1 ( .OUT(na3671_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3671_6 ( .RAM_O1(na3671_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3671_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y32     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3672_4 ( .OUT(na3672_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3672_6 ( .RAM_O2(na3672_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3672_2), .COMP_OUT(1'b0) );
// C_MX2b////      x15y41     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3673_1 ( .OUT(na3673_1), .IN1(1'b1), .IN2(~na122_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na131_1), .IN6(~na4541_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x35y48     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3674_4 ( .OUT(na3674_2), .IN1(na2600_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na197_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y47     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3675_1 ( .OUT(na3675_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2600_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na197_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x33y47     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3676_1 ( .OUT(na3676_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na4123_2), .IN7(1'b1), .IN8(na2602_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x36y47     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3677_1 ( .OUT(na3677_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na4123_2), .IN7(1'b1), .IN8(na2602_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x25y49     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3678_4 ( .OUT(na3678_2), .IN1(1'b1), .IN2(na2604_1), .IN3(1'b1), .IN4(~na197_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x27y45     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3679_1 ( .OUT(na3679_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na2604_2), .IN7(1'b1), .IN8(~na197_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x25y49     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3680_1 ( .OUT(na3680_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na951_2), .IN8(~na197_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x31y32     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3681_1 ( .OUT(na3681_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3681_6 ( .RAM_O1(na3681_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3681_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x24y62     80'h00_0018_00_0000_0888_7A5A
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3682_1 ( .OUT(na3682_1), .IN1(na3689_1), .IN2(1'b0), .IN3(~na952_1), .IN4(1'b0), .IN5(na3689_2), .IN6(1'b0), .IN7(~na952_2),
                      .IN8(~na3693_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x23y55     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3683_1 ( .OUT(na3683_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na953_2), .IN7(~na1491_1), .IN8(na864_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x31y31     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3684_4 ( .OUT(na3684_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3684_6 ( .RAM_O2(na3684_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3684_2), .COMP_OUT(1'b0) );
// C_AND////      x31y31     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3685_1 ( .OUT(na3685_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3685_6 ( .RAM_O1(na3685_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3685_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x31y30     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3686_4 ( .OUT(na3686_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3686_6 ( .RAM_O2(na3686_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3686_2), .COMP_OUT(1'b0) );
// C_AND////      x31y30     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3687_1 ( .OUT(na3687_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3687_6 ( .RAM_O1(na3687_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3687_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x37y49     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3688_4 ( .OUT(na3688_2), .IN1(1'b1), .IN2(na1593_2), .IN3(~na4523_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x23y61     80'h00_0078_00_0000_0CEE_A7B7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3689_1 ( .OUT(na3689_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na964_1), .IN6(~na2474_2), .IN7(na952_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3689_4 ( .OUT(na3689_2), .IN1(~na877_2), .IN2(~na2474_1), .IN3(na4523_2), .IN4(~na884_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y24     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3690_4 ( .OUT(na3690_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3690_6 ( .RAM_O2(na3690_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3690_2), .COMP_OUT(1'b0) );
// C_AND////      x29y24     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3691_1 ( .OUT(na3691_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3691_6 ( .RAM_O1(na3691_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3691_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///AND/      x29y23     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3692_4 ( .OUT(na3692_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3692_6 ( .RAM_O2(na3692_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3692_2), .COMP_OUT(1'b0) );
// C_MX2b////      x20y54     80'h00_0018_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3693_1 ( .OUT(na3693_1), .IN1(1'b1), .IN2(na963_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1485_1), .IN8(na2499_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x23y51     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3694_4 ( .OUT(na3694_2), .IN1(1'b1), .IN2(1'b1), .IN3(na951_1), .IN4(~na197_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x26y72     80'h00_0018_00_0000_0EEE_3557
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3695_1 ( .OUT(na3695_1), .IN1(~na1302_1), .IN2(~na929_1), .IN3(~na928_1), .IN4(1'b0), .IN5(~na1301_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(~na926_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y23     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3696_1 ( .OUT(na3696_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3696_6 ( .RAM_O1(na3696_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3696_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_///OR/      x33y72     80'h00_0060_00_0000_0C0E_FF07
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3697_4 ( .OUT(na3697_2), .IN1(~na3195_1), .IN2(~na137_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x39y71     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3698_1 ( .OUT(na3698_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na984_1), .IN6(1'b1), .IN7(na139_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x31y24     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3699_4 ( .OUT(na3699_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3699_6 ( .RAM_O2(na3699_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3699_2), .COMP_OUT(1'b0) );
// C_AND////      x13y85     80'h00_0018_00_0000_0888_2121
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3700_1 ( .OUT(na3700_1), .IN1(~na418_1), .IN2(~na412_1), .IN3(na4157_2), .IN4(~na413_1), .IN5(~na411_1), .IN6(~na4413_2),
                      .IN7(na992_1), .IN8(~na1350_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x35y82     80'h00_0060_00_0000_0C08_FF37
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3701_4 ( .OUT(na3701_2), .IN1(~na2714_1), .IN2(~na232_2), .IN3(1'b0), .IN4(~na1039_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x31y24     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3702_1 ( .OUT(na3702_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3702_6 ( .RAM_O1(na3702_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3702_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_AND////      x44y91     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3703_1 ( .OUT(na3703_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2706_1), .IN7(1'b1), .IN8(~na2707_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x31y23     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3704_4 ( .OUT(na3704_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3704_6 ( .RAM_O2(na3704_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3704_2), .COMP_OUT(1'b0) );
// C_AND////      x31y23     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3705_1 ( .OUT(na3705_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3705_6 ( .RAM_O1(na3705_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3705_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ORAND////      x42y85     80'h00_0018_00_0000_0C88_DCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3706_1 ( .OUT(na3706_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na4551_2), .IN7(~na2713_2), .IN8(na2710_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x38y82     80'h00_0018_00_0000_0C88_2FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3707_1 ( .OUT(na3707_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na2713_2), .IN8(~na2710_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x38y85     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3708_4 ( .OUT(na3708_2), .IN1(1'b0), .IN2(na1047_1), .IN3(1'b0), .IN4(na1512_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x31y22     80'h08_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3709_4 ( .OUT(na3709_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3709_6 ( .RAM_O2(na3709_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na3709_2), .COMP_OUT(1'b0) );
// C_AND////      x31y22     80'h04_0018_00_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3710_1 ( .OUT(na3710_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a3710_6 ( .RAM_O1(na3710_9), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na3710_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_////RAM_I2      x34y28     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3711_5 ( .OUT(na3711_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_93), .CP_O(1'b0) );
// C_/RAM_I1///      x34y28     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3712_2 ( .OUT(na3712_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_94), .CP_O(1'b0) );
// C_////RAM_I2      x34y27     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3713_5 ( .OUT(na3713_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_95), .CP_O(1'b0) );
// C_/RAM_I1///      x34y27     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3714_2 ( .OUT(na3714_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_96), .CP_O(1'b0) );
// C_////RAM_I2      x34y26     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3715_5 ( .OUT(na3715_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_97), .CP_O(1'b0) );
// C_/RAM_I1///      x34y26     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3716_2 ( .OUT(na3716_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_98), .CP_O(1'b0) );
// C_////RAM_I2      x34y25     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3717_5 ( .OUT(na3717_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_99), .CP_O(1'b0) );
// C_/RAM_I1///      x34y25     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3718_2 ( .OUT(na3718_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_100), .CP_O(1'b0) );
// C_////RAM_I2      x34y20     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3719_5 ( .OUT(na3719_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_113), .CP_O(1'b0) );
// C_/RAM_I1///      x34y20     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3720_2 ( .OUT(na3720_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_114), .CP_O(1'b0) );
// C_////RAM_I2      x34y19     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3721_5 ( .OUT(na3721_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_115), .CP_O(1'b0) );
// C_/RAM_I1///      x34y19     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3722_2 ( .OUT(na3722_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_116), .CP_O(1'b0) );
// C_////RAM_I2      x34y18     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3723_5 ( .OUT(na3723_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_117), .CP_O(1'b0) );
// C_/RAM_I1///      x34y18     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3724_2 ( .OUT(na3724_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_118), .CP_O(1'b0) );
// C_////RAM_I2      x34y17     80'h02_0000_00_0000_0C00_FFFF
C_RAM_I2   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3725_5 ( .OUT(na3725_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_119), .CP_O(1'b0) );
// C_/RAM_I1///      x34y17     80'h01_0000_00_0000_0C00_FFFF
C_RAM_I1   #(.CPE_CFG (9'bX_1000_0000)) 
           _a3726_2 ( .OUT(na3726_1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(na3226_120), .CP_O(1'b0) );
// C_///AND/      x45y90     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3775_4 ( .OUT(na3775_2), .IN1(na434_2), .IN2(~na2706_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x63y80     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3777_4 ( .OUT(na3777_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na38_2), .IN4(na1085_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x65y72     80'h00_0018_00_0000_0C66_C300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3778_1 ( .OUT(na3778_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1087_1), .IN7(1'b0), .IN8(na1985_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x40y69     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3782_1 ( .OUT(na3782_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na821_1), .IN6(~na817_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y71     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3783_1 ( .OUT(na3783_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4136_2), .IN5(~na1294_1), .IN6(1'b0), .IN7(~na2741_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x31y69     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3786_1 ( .OUT(na3786_1), .IN1(1'b1), .IN2(na219_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na4559_2), .IN6(~na1338_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x35y69     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3789_1 ( .OUT(na3789_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na4136_2), .IN5(~na1295_1), .IN6(1'b0), .IN7(~na2743_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y69     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3792_1 ( .OUT(na3792_1), .IN1(1'b1), .IN2(na219_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na4560_2), .IN6(~na1298_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x33y67     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3795_1 ( .OUT(na3795_1), .IN1(1'b1), .IN2(~na219_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1308_1), .IN6(~na2745_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x51y84     80'h00_0018_00_0000_0C88_A5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3796_1 ( .OUT(na3796_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na821_1), .IN6(1'b1), .IN7(na2847_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x58y82     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3797_4 ( .OUT(na3797_2), .IN1(~na821_1), .IN2(1'b1), .IN3(na2847_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y81     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3798_4 ( .OUT(na3798_2), .IN1(~na821_1), .IN2(1'b1), .IN3(na2849_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x59y85     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3799_4 ( .OUT(na3799_2), .IN1(~na821_1), .IN2(1'b1), .IN3(na2849_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x49y83     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3800_1 ( .OUT(na3800_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na821_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2851_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x47y83     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3801_1 ( .OUT(na3801_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na821_1), .IN6(1'b1), .IN7(1'b1), .IN8(na2851_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y85     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3802_1 ( .OUT(na3802_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na821_1), .IN6(na1112_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x42y92     80'h00_0018_00_0000_0888_7A3A
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3804_1 ( .OUT(na3804_1), .IN1(na3817_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na1113_1), .IN5(na3817_2), .IN6(1'b0), .IN7(~na3821_1),
                      .IN8(~na1113_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x39y85     80'h00_0060_00_0000_0C06_FFC9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3805_4 ( .OUT(na3805_2), .IN1(na1114_1), .IN2(~na1513_1), .IN3(1'b0), .IN4(na993_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x33y89     80'h00_0018_00_0000_0C66_5600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3809_1 ( .OUT(na3809_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1120_2), .IN6(na1505_2), .IN7(~na1122_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x38y87     80'h00_0060_00_0000_0C08_FF55
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3811_4 ( .OUT(na3811_2), .IN1(~na2712_1), .IN2(1'b1), .IN3(~na2713_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x33y87     80'h00_0018_00_0000_0888_AF3E
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3812_1 ( .OUT(na3812_1), .IN1(na434_1), .IN2(na4626_2), .IN3(1'b0), .IN4(~na4612_2), .IN5(1'b1), .IN6(1'b1), .IN7(na3815_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x34y87     80'h00_0078_00_0000_0C88_AA58
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3815_1 ( .OUT(na3815_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na434_2), .IN6(1'b1), .IN7(na432_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3815_4 ( .OUT(na3815_2), .IN1(na2712_2), .IN2(na4553_2), .IN3(~na2713_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x59y81     80'h00_0060_00_0000_0C08_FF2F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3816_4 ( .OUT(na3816_2), .IN1(1'b1), .IN2(1'b1), .IN3(na1599_2), .IN4(~na2707_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x39y91     80'h00_0078_00_0000_0CEE_D5B7
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3817_1 ( .OUT(na3817_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1134_1), .IN6(1'b0), .IN7(~na4548_2), .IN8(na1113_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3817_4 ( .OUT(na3817_2), .IN1(~na1037_2), .IN2(~na1047_1), .IN3(na4548_2), .IN4(~na2707_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x40y91     80'h00_0018_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3821_1 ( .OUT(na3821_1), .IN1(na1133_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1507_1), .IN8(na2739_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x51y84     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3822_4 ( .OUT(na3822_2), .IN1(~na821_1), .IN2(na1112_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x49y76     80'h00_0018_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3823_1 ( .OUT(na3823_1), .IN1(1'b1), .IN2(~na285_1), .IN3(1'b0), .IN4(1'b0), .IN5(na21_1), .IN6(na3159_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x58y83     80'h00_0018_00_0000_0C88_BCFF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3826_1 ( .OUT(na3826_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(na2965_2), .IN7(na2961_1), .IN8(~na4571_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x59y83     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3827_1 ( .OUT(na3827_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na2962_2), .IN6(1'b1), .IN7(~na2961_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x65y87     80'h00_0018_00_0000_0C66_6000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3828_1 ( .OUT(na3828_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1534_2), .IN8(na1195_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x61y87     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3895_1 ( .OUT(na3895_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na2957_2), .IN6(1'b1), .IN7(1'b1), .IN8(na986_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x20y61     80'h00_0060_00_0000_0C08_FF53
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3898_4 ( .OUT(na3898_2), .IN1(1'b1), .IN2(~na421_1), .IN3(~na426_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x21y65     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3899_1 ( .OUT(na3899_1), .IN1(1'b1), .IN2(na423_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2986_1), .IN6(~na1320_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x21y67     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3902_1 ( .OUT(na3902_1), .IN1(1'b1), .IN2(na423_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2986_2), .IN6(~na633_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x25y63     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3905_1 ( .OUT(na3905_1), .IN1(1'b1), .IN2(~na423_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na634_1), .IN6(~na4578_2), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x19y65     80'h00_0018_00_0040_0A33_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3908_1 ( .OUT(na3908_1), .IN1(1'b1), .IN2(na423_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na2988_2), .IN6(~na635_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x17y65     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3911_1 ( .OUT(na3911_1), .IN1(1'b1), .IN2(~na423_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na1319_1), .IN6(~na2990_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x33y63     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3912_4 ( .OUT(na3912_2), .IN1(na3105_1), .IN2(1'b1), .IN3(~na426_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x35y63     80'h00_0060_00_0000_0C08_FF5A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3913_4 ( .OUT(na3913_2), .IN1(na3105_2), .IN2(1'b1), .IN3(~na426_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x33y63     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3914_1 ( .OUT(na3914_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3107_1), .IN6(1'b1), .IN7(~na426_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y63     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3915_1 ( .OUT(na3915_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na3107_2), .IN6(1'b1), .IN7(~na426_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y62     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3916_1 ( .OUT(na3916_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na426_1), .IN8(na3109_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x39y61     80'h00_0060_00_0000_0C08_FF4F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3917_4 ( .OUT(na3917_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na426_1), .IN4(na3109_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x42y66     80'h00_0060_00_0000_0C08_FF5C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3918_4 ( .OUT(na3918_2), .IN1(1'b1), .IN2(na1254_2), .IN3(~na426_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x64y85     80'h00_0018_00_0000_0888_C7C5
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3920_1 ( .OUT(na3920_1), .IN1(~na1255_1), .IN2(1'b0), .IN3(1'b0), .IN4(na3933_1), .IN5(~na1255_2), .IN6(~na3937_1), .IN7(1'b0),
                      .IN8(na3933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x64y80     80'h00_0060_00_0000_0C06_FFC9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3921_4 ( .OUT(na3921_2), .IN1(~na1535_1), .IN2(na1256_2), .IN3(1'b0), .IN4(na1388_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x50y88     80'h00_0018_00_0000_0C66_6300
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3925_1 ( .OUT(na3925_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1264_1), .IN7(na1527_2), .IN8(na1262_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x61y83     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3927_4 ( .OUT(na3927_2), .IN1(~na2963_2), .IN2(~na2965_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x57y90     80'h00_0018_00_0000_0888_FAE3
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a3928_1 ( .OUT(na3928_1), .IN1(1'b0), .IN2(~na4589_2), .IN3(na4629_2), .IN4(na986_1), .IN5(na3931_2), .IN6(1'b0), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x55y87     80'h00_0078_00_0000_0C88_8FC2
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3931_1 ( .OUT(na3931_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na980_2), .IN8(na986_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3931_4 ( .OUT(na3931_2), .IN1(na2962_1), .IN2(~na2965_2), .IN3(1'b1), .IN4(na4571_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x55y82     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3932_1 ( .OUT(na3932_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2958_2), .IN8(na1605_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x66y86     80'h00_0078_00_0000_0CEE_7A7D
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3933_1 ( .OUT(na3933_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1255_2), .IN6(1'b0), .IN7(~na2958_2), .IN8(~na1276_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a3933_4 ( .OUT(na3933_2), .IN1(~na460_2), .IN2(na4566_2), .IN3(~na2958_1), .IN4(~na1195_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x59y88     80'h00_0018_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3937_1 ( .OUT(na3937_1), .IN1(1'b1), .IN2(~na1275_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na2984_1), .IN8(na1529_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x39y67     80'h00_0018_00_0000_0C88_5CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3938_1 ( .OUT(na3938_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1254_1), .IN7(~na426_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x25y72     80'h00_0018_00_0000_0CEE_5300
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3939_1 ( .OUT(na3939_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na3217_1), .IN7(~na4109_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x39y71     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3940_4 ( .OUT(na3940_2), .IN1(na1290_1), .IN2(1'b1), .IN3(na139_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x37y78     80'h00_0078_00_0000_0C88_3A8C
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3943_1 ( .OUT(na3943_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1188_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1296_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3943_4 ( .OUT(na3943_2), .IN1(1'b1), .IN2(na3823_1), .IN3(na506_2), .IN4(na1296_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x31y73     80'h00_0060_00_0000_0C08_FF75
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a3944_4 ( .OUT(na3944_2), .IN1(~na1188_1), .IN2(1'b0), .IN3(~na4632_2), .IN4(~na1296_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x49y67     80'h00_0018_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3948_1 ( .OUT(na3948_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1314_2), .IN6(1'b1), .IN7(na139_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x24y67     80'h00_0060_00_0000_0C08_FFA3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3950_4 ( .OUT(na3950_2), .IN1(1'b1), .IN2(~na405_2), .IN3(na233_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x33y81     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3954_1 ( .OUT(na3954_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na232_2), .IN7(1'b1), .IN8(na1341_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x47y88     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3955_4 ( .OUT(na3955_2), .IN1(~na1343_1), .IN2(na2706_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x26y84     80'h00_0018_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3958_1 ( .OUT(na3958_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na287_2), .IN8(na1296_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y66     80'h00_0060_00_0000_0C08_FF3A
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3960_4 ( .OUT(na3960_2), .IN1(na1370_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na214_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x23y59     80'h00_0060_00_0000_0C06_FFC5
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3961_4 ( .OUT(na3961_2), .IN1(~na1372_1), .IN2(1'b0), .IN3(1'b0), .IN4(na2473_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x48y61     80'h00_0018_00_0000_0EEE_3077
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a3964_1 ( .OUT(na3964_1), .IN1(~na1387_1), .IN2(~na1386_1), .IN3(~na283_1), .IN4(~na284_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                      .IN8(~na282_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x51y59     80'h00_0018_00_0000_0888_1555
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3975_1 ( .OUT(na3975_1), .IN1(~na2001_2), .IN2(1'b1), .IN3(~na2002_1), .IN4(1'b1), .IN5(~na2001_1), .IN6(1'b1), .IN7(~na1999_1),
                      .IN8(~na2000_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x69y74     80'h00_0018_00_0040_0C86_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3977_1 ( .OUT(na3977_1), .IN1(1'b0), .IN2(na1438_1), .IN3(na4420_2), .IN4(1'b1), .IN5(na524_1), .IN6(1'b1), .IN7(na520_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x67y80     80'h00_0018_00_0040_0C86_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3978_1 ( .OUT(na3978_1), .IN1(1'b0), .IN2(na4421_2), .IN3(na1439_1), .IN4(1'b1), .IN5(~na607_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na605_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x55y86     80'h00_0018_00_0040_0C49_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3979_1 ( .OUT(na3979_1), .IN1(na4422_2), .IN2(1'b0), .IN3(1'b1), .IN4(na1440_2), .IN5(~na4080_2), .IN6(1'b1), .IN7(na613_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x65y65     80'h00_0018_00_0040_0A68_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3981_1 ( .OUT(na3981_1), .IN1(1'b1), .IN2(~na599_2), .IN3(na4226_2), .IN4(1'b1), .IN5(1'b0), .IN6(na4427_2), .IN7(na1447_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x68y65     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3983_1 ( .OUT(na3983_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2350_2), .IN7(1'b1), .IN8(~na1985_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x52y46     80'h00_0018_00_0000_0888_3313
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a3988_1 ( .OUT(na3988_1), .IN1(1'b1), .IN2(~na2238_1), .IN3(~na2239_1), .IN4(~na2237_2), .IN5(1'b1), .IN6(~na2238_2), .IN7(1'b1),
                      .IN8(~na2236_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x61y59     80'h00_0018_00_0040_0C49_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3990_1 ( .OUT(na3990_1), .IN1(na4429_2), .IN2(1'b0), .IN3(1'b1), .IN4(na1460_2), .IN5(~na708_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na4262_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x61y70     80'h00_0018_00_0040_0C49_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3991_1 ( .OUT(na3991_1), .IN1(na4430_2), .IN2(1'b0), .IN3(1'b1), .IN4(na1461_1), .IN5(na253_1), .IN6(1'b1), .IN7(na251_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x53y73     80'h00_0018_00_0040_0C86_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3992_1 ( .OUT(na3992_1), .IN1(1'b0), .IN2(na4431_2), .IN3(na1462_2), .IN4(1'b1), .IN5(1'b1), .IN6(na261_2), .IN7(1'b1), .IN8(na327_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y50     80'h00_0018_00_0040_0A68_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a3994_1 ( .OUT(na3994_1), .IN1(1'b1), .IN2(~na786_1), .IN3(1'b1), .IN4(na720_1), .IN5(1'b0), .IN6(na4436_2), .IN7(na1469_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x65y47     80'h00_0060_00_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a3996_4 ( .OUT(na3996_2), .IN1(~na704_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na4503_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x20y40     80'h00_0018_00_0000_0888_1F15
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4001_1 ( .OUT(na4001_1), .IN1(~na2490_2), .IN2(1'b1), .IN3(~na2488_1), .IN4(~na2489_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na2487_2),
                      .IN8(~na2489_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x18y57     80'h00_0018_00_0040_0C86_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4003_1 ( .OUT(na4003_1), .IN1(1'b0), .IN2(na1482_2), .IN3(na4438_2), .IN4(1'b1), .IN5(na882_2), .IN6(1'b1), .IN7(1'b1), .IN8(na885_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x19y66     80'h00_0018_00_0040_0C49_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4004_1 ( .OUT(na4004_1), .IN1(na1483_2), .IN2(1'b0), .IN3(1'b1), .IN4(na4439_2), .IN5(1'b1), .IN6(na180_1), .IN7(1'b1), .IN8(na178_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x15y72     80'h00_0018_00_0040_0C49_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4005_1 ( .OUT(na4005_1), .IN1(na1484_2), .IN2(1'b0), .IN3(1'b1), .IN4(na4440_2), .IN5(1'b1), .IN6(~na119_1), .IN7(1'b1),
                      .IN8(na188_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x22y56     80'h00_0018_00_0040_0A68_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4007_1 ( .OUT(na4007_1), .IN1(1'b1), .IN2(~na953_2), .IN3(1'b1), .IN4(na864_1), .IN5(1'b0), .IN6(na4446_2), .IN7(na1491_1),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x34y49     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4009_1 ( .OUT(na4009_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na881_2), .IN7(1'b1), .IN8(~na2473_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x38y70     80'h00_0018_00_0000_0888_1535
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4014_1 ( .OUT(na4014_1), .IN1(~na4556_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na2722_1), .IN5(~na4555_2), .IN6(1'b1), .IN7(~na4557_2),
                      .IN8(~na2723_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x40y90     80'h00_0018_00_0040_0C86_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4016_1 ( .OUT(na4016_1), .IN1(1'b0), .IN2(na1504_2), .IN3(na4447_2), .IN4(1'b1), .IN5(na1045_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na1049_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x31y91     80'h00_0018_00_0040_0C86_5A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4017_1 ( .OUT(na4017_1), .IN1(1'b0), .IN2(na1505_2), .IN3(na4448_2), .IN4(1'b1), .IN5(na1120_2), .IN6(1'b1), .IN7(~na1122_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x27y91     80'h00_0018_00_0040_0C16_3500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4018_1 ( .OUT(na4018_1), .IN1(1'b1), .IN2(na1506_1), .IN3(na4449_2), .IN4(1'b0), .IN5(~na1292_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na1128_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x35y83     80'h00_0018_00_0040_0A68_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4020_1 ( .OUT(na4020_1), .IN1(~na1114_1), .IN2(1'b1), .IN3(1'b1), .IN4(na993_1), .IN5(1'b0), .IN6(na1513_1), .IN7(na4452_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x57y86     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4022_4 ( .OUT(na4022_2), .IN1(1'b1), .IN2(~na1044_2), .IN3(1'b1), .IN4(~na4544_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x31y66     80'h00_0018_00_0000_0888_3351
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4027_1 ( .OUT(na4027_1), .IN1(~na2974_2), .IN2(~na2973_2), .IN3(~na2972_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na2973_1), .IN7(1'b1),
                      .IN8(~na2971_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x63y88     80'h00_0018_00_0040_0C49_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4029_1 ( .OUT(na4029_1), .IN1(na4453_2), .IN2(1'b0), .IN3(1'b1), .IN4(na1526_1), .IN5(~na1197_1), .IN6(1'b1), .IN7(na4370_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x49y91     80'h00_0018_00_0040_0C86_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4030_1 ( .OUT(na4030_1), .IN1(1'b0), .IN2(na4454_2), .IN3(na1527_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na1264_1), .IN7(1'b1),
                      .IN8(na1262_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x48y91     80'h00_0018_00_0040_0C86_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4031_1 ( .OUT(na4031_1), .IN1(1'b0), .IN2(na1528_2), .IN3(na4455_2), .IN4(1'b1), .IN5(na1270_2), .IN6(1'b1), .IN7(1'b1),
                      .IN8(na532_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x61y80     80'h00_0018_00_0040_0A94_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a4033_1 ( .OUT(na4033_1), .IN1(1'b1), .IN2(na1256_2), .IN3(1'b1), .IN4(na1388_1), .IN5(na1535_1), .IN6(1'b0), .IN7(1'b1),
                      .IN8(na4459_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x67y81     80'h00_0060_00_0000_0C08_FFF1
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4035_4 ( .OUT(na4035_2), .IN1(~na1192_2), .IN2(~na4563_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x68y81     80'h00_0078_00_0000_0C66_3ACC
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4039_1 ( .OUT(na4039_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2091_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na76_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4039_4 ( .OUT(na4039_2), .IN1(1'b0), .IN2(na2093_1), .IN3(1'b0), .IN4(na76_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x67y83     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4040_1 ( .OUT(na4040_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2091_2), .IN6(~na75_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x65y81     80'h00_0018_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4041_1 ( .OUT(na4041_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na534_2), .IN6(1'b1), .IN7(1'b1), .IN8(na78_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x70y82     80'h00_0060_00_0000_0C06_FFCA
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4042_4 ( .OUT(na4042_2), .IN1(na534_1), .IN2(1'b0), .IN3(1'b0), .IN4(na78_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x71y79     80'h00_0018_00_0000_0EEE_ED7B
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a4043_1 ( .OUT(na4043_1), .IN1(na4041_1), .IN2(~na94_1), .IN3(~na4039_1), .IN4(~na50_1), .IN5(~na4040_1), .IN6(na94_2), .IN7(na4039_2),
                      .IN8(na4042_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x17y87     80'h00_0078_00_0000_0C66_095A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4045_1 ( .OUT(na4045_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na390_2), .IN6(na1051_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4045_4 ( .OUT(na4045_2), .IN1(na2819_1), .IN2(1'b0), .IN3(~na388_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x22y91     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4046_1 ( .OUT(na4046_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na390_1), .IN6(na1051_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x16y53     80'h00_0078_00_0000_0C66_A5A5
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4050_1 ( .OUT(na4050_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na192_2), .IN6(1'b0), .IN7(na891_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4050_4 ( .OUT(na4050_2), .IN1(~na192_1), .IN2(1'b0), .IN3(na891_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x37y60     80'h00_0078_00_0000_0C66_90C3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4053_1 ( .OUT(na4053_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na264_1), .IN8(na2337_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4053_4 ( .OUT(na4053_2), .IN1(1'b0), .IN2(~na265_2), .IN3(1'b0), .IN4(na2337_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x48y53     80'h00_0060_00_0000_0C06_FFA3
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4054_4 ( .OUT(na4054_2), .IN1(1'b0), .IN2(~na265_1), .IN3(na2339_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x63y92     80'h00_0078_00_0000_0C66_A390
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4058_1 ( .OUT(na4058_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na825_1), .IN7(na3064_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4058_4 ( .OUT(na4058_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3064_1), .IN4(~na826_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x68y91     80'h00_0060_00_0000_0C06_FF3C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4059_4 ( .OUT(na4059_2), .IN1(1'b0), .IN2(na3066_1), .IN3(1'b0), .IN4(~na826_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x15y47     80'h00_0078_00_0000_0C66_A590
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4063_1 ( .OUT(na4063_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na173_1), .IN6(1'b0), .IN7(na2579_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4063_4 ( .OUT(na4063_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2579_1), .IN4(~na190_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x15y52     80'h00_0018_00_0000_0C66_9000
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4064_1 ( .OUT(na4064_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na4120_2), .IN8(na2581_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x1y51     80'h08_0060_00_0000_0C08_FFF5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a4065_4 ( .OUT(na4065_2), .IN1(~na1540_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a4065_6 ( .RAM_O2(na4065_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na4065_2), .COMP_OUT(1'b0) );
// C_////Bridge      x52y70     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4066_5 ( .OUT(na4066_2), .IN1(1'b0), .IN2(na12_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4067_5 ( .OUT(na4067_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na16_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4068_5 ( .OUT(na4068_2), .IN1(1'b0), .IN2(1'b0), .IN3(na17_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y48     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4069_5 ( .OUT(na4069_2), .IN1(1'b0), .IN2(1'b0), .IN3(na17_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4070_5 ( .OUT(na4070_2), .IN1(1'b0), .IN2(na22_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y68     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4071_5 ( .OUT(na4071_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na27_1) );
// C_////Bridge      x21y70     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4072_5 ( .OUT(na4072_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na27_2) );
// C_////Bridge      x24y65     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4073_5 ( .OUT(na4073_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na28_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y79     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4074_5 ( .OUT(na4074_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na30_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y62     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4075_5 ( .OUT(na4075_2), .IN1(na31_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y70     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4076_5 ( .OUT(na4076_2), .IN1(1'b0), .IN2(na33_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y71     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4077_5 ( .OUT(na4077_2), .IN1(1'b0), .IN2(1'b0), .IN3(na38_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y77     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4078_5 ( .OUT(na4078_2), .IN1(1'b0), .IN2(1'b0), .IN3(na38_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y75     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4079_5 ( .OUT(na4079_2), .IN1(1'b0), .IN2(na40_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y85     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4080_5 ( .OUT(na4080_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na46_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y85     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4081_5 ( .OUT(na4081_2), .IN1(1'b0), .IN2(na47_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y75     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4082_5 ( .OUT(na4082_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na51_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y75     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4083_5 ( .OUT(na4083_2), .IN1(na53_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y57     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4084_5 ( .OUT(na4084_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na54_2) );
// C_////Bridge      x61y81     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4085_5 ( .OUT(na4085_2), .IN1(1'b0), .IN2(na57_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y83     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4086_5 ( .OUT(na4086_2), .IN1(1'b0), .IN2(na58_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y75     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4087_5 ( .OUT(na4087_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na67_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y71     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4088_5 ( .OUT(na4088_2), .IN1(1'b0), .IN2(1'b0), .IN3(na70_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4089_5 ( .OUT(na4089_2), .IN1(1'b0), .IN2(1'b0), .IN3(na85_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4090_5 ( .OUT(na4090_2), .IN1(na90_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y50     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4091_5 ( .OUT(na4091_2), .IN1(1'b0), .IN2(na91_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y50     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4092_5 ( .OUT(na4092_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na93_1), .IN8(1'b0) );
// C_////Bridge      x38y55     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4093_5 ( .OUT(na4093_2), .IN1(1'b0), .IN2(na94_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4094_5 ( .OUT(na4094_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na104_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y75     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4095_5 ( .OUT(na4095_2), .IN1(1'b0), .IN2(1'b0), .IN3(na107_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y54     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4096_5 ( .OUT(na4096_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na108_1) );
// C_////Bridge      x62y75     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4097_5 ( .OUT(na4097_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na109_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y65     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4098_5 ( .OUT(na4098_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na110_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4099_5 ( .OUT(na4099_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na112_1) );
// C_////Bridge      x18y62     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4100_5 ( .OUT(na4100_2), .IN1(na114_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y75     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4101_5 ( .OUT(na4101_2), .IN1(1'b0), .IN2(1'b0), .IN3(na115_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4102_5 ( .OUT(na4102_2), .IN1(1'b0), .IN2(1'b0), .IN3(na115_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4103_5 ( .OUT(na4103_2), .IN1(na117_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x14y69     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4104_5 ( .OUT(na4104_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na120_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y57     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4105_5 ( .OUT(na4105_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na124_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4106_5 ( .OUT(na4106_2), .IN1(na129_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y75     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4107_5 ( .OUT(na4107_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na133_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y84     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4108_5 ( .OUT(na4108_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na135_1) );
// C_////Bridge      x30y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4109_5 ( .OUT(na4109_2), .IN1(1'b0), .IN2(na137_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y79     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4110_5 ( .OUT(na4110_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na139_1), .IN8(1'b0) );
// C_////Bridge      x60y68     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4111_5 ( .OUT(na4111_2), .IN1(na145_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y85     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4112_5 ( .OUT(na4112_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na158_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y83     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4113_5 ( .OUT(na4113_2), .IN1(na160_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x15y82     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4114_5 ( .OUT(na4114_2), .IN1(na163_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4115_5 ( .OUT(na4115_2), .IN1(na166_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4116_5 ( .OUT(na4116_2), .IN1(na167_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4117_5 ( .OUT(na4117_2), .IN1(na169_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y79     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4118_5 ( .OUT(na4118_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na170_1) );
// C_////Bridge      x15y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4119_5 ( .OUT(na4119_2), .IN1(1'b0), .IN2(1'b0), .IN3(na189_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x16y51     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4120_5 ( .OUT(na4120_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na190_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x16y48     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4121_5 ( .OUT(na4121_2), .IN1(1'b0), .IN2(na193_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y42     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4122_5 ( .OUT(na4122_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na194_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y46     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4123_5 ( .OUT(na4123_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na197_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y38     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4124_5 ( .OUT(na4124_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na203_1) );
// C_////Bridge      x27y45     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4125_5 ( .OUT(na4125_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na203_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y39     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4126_5 ( .OUT(na4126_2), .IN1(1'b0), .IN2(na207_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y37     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4127_5 ( .OUT(na4127_2), .IN1(1'b0), .IN2(na207_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4128_5 ( .OUT(na4128_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na208_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x15y59     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4129_5 ( .OUT(na4129_2), .IN1(1'b0), .IN2(na209_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y54     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4130_5 ( .OUT(na4130_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na211_1), .IN8(1'b0) );
// C_////Bridge      x21y61     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4131_5 ( .OUT(na4131_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na214_1) );
// C_////Bridge      x27y54     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4132_5 ( .OUT(na4132_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na214_2) );
// C_////Bridge      x36y51     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4133_5 ( .OUT(na4133_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na216_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x18y59     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4134_5 ( .OUT(na4134_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na216_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4135_5 ( .OUT(na4135_2), .IN1(na218_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y70     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4136_5 ( .OUT(na4136_2), .IN1(1'b0), .IN2(na219_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4137_5 ( .OUT(na4137_2), .IN1(na220_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4138_5 ( .OUT(na4138_2), .IN1(na222_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y90     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4139_5 ( .OUT(na4139_2), .IN1(1'b0), .IN2(na225_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y77     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4140_5 ( .OUT(na4140_2), .IN1(1'b0), .IN2(na232_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y81     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4141_5 ( .OUT(na4141_2), .IN1(1'b0), .IN2(na232_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4142_5 ( .OUT(na4142_2), .IN1(1'b0), .IN2(1'b0), .IN3(na233_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x13y66     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4143_5 ( .OUT(na4143_2), .IN1(1'b0), .IN2(1'b0), .IN3(na233_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y80     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4144_5 ( .OUT(na4144_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na240_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y87     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4145_5 ( .OUT(na4145_2), .IN1(1'b0), .IN2(1'b0), .IN3(na241_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4146_5 ( .OUT(na4146_2), .IN1(na243_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y71     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4147_5 ( .OUT(na4147_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na245_1) );
// C_////Bridge      x61y77     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4148_5 ( .OUT(na4148_2), .IN1(1'b0), .IN2(1'b0), .IN3(na246_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y33     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4149_5 ( .OUT(na4149_2), .IN1(1'b0), .IN2(1'b0), .IN3(na280_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y35     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4150_5 ( .OUT(na4150_2), .IN1(1'b0), .IN2(1'b0), .IN3(na280_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4151_5 ( .OUT(na4151_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na282_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4152_5 ( .OUT(na4152_2), .IN1(1'b0), .IN2(na285_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y68     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4153_5 ( .OUT(na4153_2), .IN1(1'b0), .IN2(na285_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y64     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4154_5 ( .OUT(na4154_2), .IN1(1'b0), .IN2(na285_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y76     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4155_5 ( .OUT(na4155_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na287_2), .IN8(1'b0) );
// C_////Bridge      x18y80     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4156_5 ( .OUT(na4156_2), .IN1(1'b0), .IN2(na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x16y85     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4157_5 ( .OUT(na4157_2), .IN1(1'b0), .IN2(na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x18y82     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4158_5 ( .OUT(na4158_2), .IN1(1'b0), .IN2(na288_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y62     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4159_5 ( .OUT(na4159_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na295_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y58     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4160_5 ( .OUT(na4160_2), .IN1(1'b0), .IN2(na295_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y55     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4161_5 ( .OUT(na4161_2), .IN1(1'b0), .IN2(1'b0), .IN3(na297_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4162_5 ( .OUT(na4162_2), .IN1(1'b0), .IN2(1'b0), .IN3(na297_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x13y61     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4163_5 ( .OUT(na4163_2), .IN1(1'b0), .IN2(na299_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y58     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4164_5 ( .OUT(na4164_2), .IN1(1'b0), .IN2(na299_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y42     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4165_5 ( .OUT(na4165_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na303_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x16y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4166_5 ( .OUT(na4166_2), .IN1(1'b0), .IN2(1'b0), .IN3(na304_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y76     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4167_5 ( .OUT(na4167_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na311_1), .IN8(1'b0) );
// C_////Bridge      x29y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4168_5 ( .OUT(na4168_2), .IN1(na316_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4169_5 ( .OUT(na4169_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na322_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y67     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4170_5 ( .OUT(na4170_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na324_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y64     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4171_5 ( .OUT(na4171_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na331_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y62     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4172_5 ( .OUT(na4172_2), .IN1(1'b0), .IN2(1'b0), .IN3(na332_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y62     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4173_5 ( .OUT(na4173_2), .IN1(na333_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y56     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4174_5 ( .OUT(na4174_2), .IN1(na335_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4175_5 ( .OUT(na4175_2), .IN1(1'b0), .IN2(1'b0), .IN3(na353_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y55     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4176_5 ( .OUT(na4176_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na354_1), .IN8(1'b0) );
// C_////Bridge      x70y54     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4177_5 ( .OUT(na4177_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na355_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y56     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4178_5 ( .OUT(na4178_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na356_1), .IN8(1'b0) );
// C_////Bridge      x26y55     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4179_5 ( .OUT(na4179_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na358_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y76     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4180_5 ( .OUT(na4180_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na360_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y77     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4181_5 ( .OUT(na4181_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na362_2), .IN8(1'b0) );
// C_////Bridge      x43y75     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4182_5 ( .OUT(na4182_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na363_2), .IN8(1'b0) );
// C_////Bridge      x35y70     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4183_5 ( .OUT(na4183_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na364_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y71     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4184_5 ( .OUT(na4184_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na365_2), .IN8(1'b0) );
// C_////Bridge      x45y74     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4185_5 ( .OUT(na4185_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na366_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y73     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4186_5 ( .OUT(na4186_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na367_2), .IN8(1'b0) );
// C_////Bridge      x45y75     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4187_5 ( .OUT(na4187_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na368_2), .IN8(1'b0) );
// C_////Bridge      x43y78     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4188_5 ( .OUT(na4188_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na369_2) );
// C_////Bridge      x26y89     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4189_5 ( .OUT(na4189_2), .IN1(na370_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y87     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4190_5 ( .OUT(na4190_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na371_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y90     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4191_5 ( .OUT(na4191_2), .IN1(na374_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y89     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4192_5 ( .OUT(na4192_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na409_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y86     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4193_5 ( .OUT(na4193_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na410_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y56     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4194_5 ( .OUT(na4194_2), .IN1(1'b0), .IN2(na421_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y72     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4195_5 ( .OUT(na4195_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na424_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y72     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4196_5 ( .OUT(na4196_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na428_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4197_5 ( .OUT(na4197_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na429_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y91     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4198_5 ( .OUT(na4198_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na432_2), .IN8(1'b0) );
// C_////Bridge      x34y93     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4199_5 ( .OUT(na4199_2), .IN1(na434_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4200_5 ( .OUT(na4200_2), .IN1(na434_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4201_5 ( .OUT(na4201_2), .IN1(1'b0), .IN2(1'b0), .IN3(na443_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4202_5 ( .OUT(na4202_2), .IN1(na445_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4203_5 ( .OUT(na4203_2), .IN1(na445_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y90     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4204_5 ( .OUT(na4204_2), .IN1(na455_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y68     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4205_5 ( .OUT(na4205_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na456_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4206_5 ( .OUT(na4206_2), .IN1(na456_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4207_5 ( .OUT(na4207_2), .IN1(na456_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y87     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4208_5 ( .OUT(na4208_2), .IN1(1'b0), .IN2(1'b0), .IN3(na461_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4209_5 ( .OUT(na4209_2), .IN1(1'b0), .IN2(1'b0), .IN3(na461_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y52     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4210_5 ( .OUT(na4210_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na465_1), .IN8(1'b0) );
// C_////Bridge      x68y85     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4211_5 ( .OUT(na4211_2), .IN1(1'b0), .IN2(na466_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y76     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4212_5 ( .OUT(na4212_2), .IN1(1'b0), .IN2(na469_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y66     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4213_5 ( .OUT(na4213_2), .IN1(na486_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y87     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4214_5 ( .OUT(na4214_2), .IN1(1'b0), .IN2(na510_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y65     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4215_5 ( .OUT(na4215_2), .IN1(1'b0), .IN2(na512_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y80     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4216_5 ( .OUT(na4216_2), .IN1(1'b0), .IN2(na512_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y72     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4217_5 ( .OUT(na4217_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na516_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x69y69     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4218_5 ( .OUT(na4218_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na517_2) );
// C_////Bridge      x66y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4219_5 ( .OUT(na4219_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na519_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y64     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4220_5 ( .OUT(na4220_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na519_2) );
// C_////Bridge      x72y75     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4221_5 ( .OUT(na4221_2), .IN1(na522_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y78     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4222_5 ( .OUT(na4222_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na523_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y50     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4223_5 ( .OUT(na4223_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na526_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y60     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4224_5 ( .OUT(na4224_2), .IN1(1'b0), .IN2(1'b0), .IN3(na529_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y85     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4225_5 ( .OUT(na4225_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na533_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y67     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4226_5 ( .OUT(na4226_2), .IN1(na535_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y38     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4227_5 ( .OUT(na4227_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na536_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y40     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4228_5 ( .OUT(na4228_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na536_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y50     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4229_5 ( .OUT(na4229_2), .IN1(na543_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y48     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4230_5 ( .OUT(na4230_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na543_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y53     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4231_5 ( .OUT(na4231_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na547_1), .IN8(1'b0) );
// C_////Bridge      x71y53     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4232_5 ( .OUT(na4232_2), .IN1(1'b0), .IN2(1'b0), .IN3(na547_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y49     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4233_5 ( .OUT(na4233_2), .IN1(1'b0), .IN2(1'b0), .IN3(na549_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y47     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4234_5 ( .OUT(na4234_2), .IN1(1'b0), .IN2(1'b0), .IN3(na549_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y49     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4235_5 ( .OUT(na4235_2), .IN1(1'b0), .IN2(1'b0), .IN3(na551_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x69y55     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4236_5 ( .OUT(na4236_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na551_2), .IN8(1'b0) );
// C_////Bridge      x65y51     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4237_5 ( .OUT(na4237_2), .IN1(1'b0), .IN2(na553_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x69y47     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4238_5 ( .OUT(na4238_2), .IN1(1'b0), .IN2(na553_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y44     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4239_5 ( .OUT(na4239_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na555_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y46     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4240_5 ( .OUT(na4240_2), .IN1(na555_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y44     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4241_5 ( .OUT(na4241_2), .IN1(na557_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y44     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4242_5 ( .OUT(na4242_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na557_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y51     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4243_5 ( .OUT(na4243_2), .IN1(1'b0), .IN2(na559_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y51     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4244_5 ( .OUT(na4244_2), .IN1(1'b0), .IN2(na559_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y49     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4245_5 ( .OUT(na4245_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na561_1), .IN8(1'b0) );
// C_////Bridge      x71y47     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4246_5 ( .OUT(na4246_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na561_2), .IN8(1'b0) );
// C_////Bridge      x66y46     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4247_5 ( .OUT(na4247_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na569_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y48     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4248_5 ( .OUT(na4248_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na569_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y46     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4249_5 ( .OUT(na4249_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na571_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y46     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4250_5 ( .OUT(na4250_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na571_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y44     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4251_5 ( .OUT(na4251_2), .IN1(na573_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y44     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4252_5 ( .OUT(na4252_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na573_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y73     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4253_5 ( .OUT(na4253_2), .IN1(1'b0), .IN2(1'b0), .IN3(na603_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y71     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4254_5 ( .OUT(na4254_2), .IN1(1'b0), .IN2(na633_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y34     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4255_5 ( .OUT(na4255_2), .IN1(1'b0), .IN2(1'b0), .IN3(na636_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4256_5 ( .OUT(na4256_2), .IN1(na647_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y59     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4257_5 ( .OUT(na4257_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na664_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y44     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4258_5 ( .OUT(na4258_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na677_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y86     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4259_5 ( .OUT(na4259_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na693_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y88     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4260_5 ( .OUT(na4260_2), .IN1(na696_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x74y43     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4261_5 ( .OUT(na4261_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na704_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y58     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4262_5 ( .OUT(na4262_2), .IN1(1'b0), .IN2(na705_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y61     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4263_5 ( .OUT(na4263_2), .IN1(na707_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y84     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4264_5 ( .OUT(na4264_2), .IN1(na712_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y45     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4265_5 ( .OUT(na4265_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na720_1) );
// C_////Bridge      x21y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4266_5 ( .OUT(na4266_2), .IN1(na727_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x73y43     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4267_5 ( .OUT(na4267_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na728_1) );
// C_////Bridge      x62y39     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4268_5 ( .OUT(na4268_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na728_2) );
// C_////Bridge      x60y43     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4269_5 ( .OUT(na4269_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na734_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y41     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4270_5 ( .OUT(na4270_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na734_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y36     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4271_5 ( .OUT(na4271_2), .IN1(1'b0), .IN2(1'b0), .IN3(na738_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y36     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4272_5 ( .OUT(na4272_2), .IN1(1'b0), .IN2(1'b0), .IN3(na738_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y38     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4273_5 ( .OUT(na4273_2), .IN1(1'b0), .IN2(1'b0), .IN3(na740_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y38     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4274_5 ( .OUT(na4274_2), .IN1(1'b0), .IN2(1'b0), .IN3(na740_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y38     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4275_5 ( .OUT(na4275_2), .IN1(1'b0), .IN2(1'b0), .IN3(na742_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y40     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4276_5 ( .OUT(na4276_2), .IN1(1'b0), .IN2(1'b0), .IN3(na742_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y38     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4277_5 ( .OUT(na4277_2), .IN1(1'b0), .IN2(1'b0), .IN3(na744_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y40     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4278_5 ( .OUT(na4278_2), .IN1(1'b0), .IN2(1'b0), .IN3(na744_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y37     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4279_5 ( .OUT(na4279_2), .IN1(1'b0), .IN2(1'b0), .IN3(na746_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y35     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4280_5 ( .OUT(na4280_2), .IN1(1'b0), .IN2(1'b0), .IN3(na746_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y39     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4281_5 ( .OUT(na4281_2), .IN1(1'b0), .IN2(1'b0), .IN3(na748_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y37     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4282_5 ( .OUT(na4282_2), .IN1(1'b0), .IN2(1'b0), .IN3(na748_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y37     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4283_5 ( .OUT(na4283_2), .IN1(na752_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y33     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4284_5 ( .OUT(na4284_2), .IN1(na752_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y33     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4285_5 ( .OUT(na4285_2), .IN1(1'b0), .IN2(na754_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y37     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4286_5 ( .OUT(na4286_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na754_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y35     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4287_5 ( .OUT(na4287_2), .IN1(1'b0), .IN2(na756_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y35     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4288_5 ( .OUT(na4288_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na756_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y38     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4289_5 ( .OUT(na4289_2), .IN1(1'b0), .IN2(1'b0), .IN3(na758_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y40     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4290_5 ( .OUT(na4290_2), .IN1(1'b0), .IN2(1'b0), .IN3(na758_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4291_5 ( .OUT(na4291_2), .IN1(na762_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y78     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4292_5 ( .OUT(na4292_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na815_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y69     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4293_5 ( .OUT(na4293_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na817_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y82     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4294_5 ( .OUT(na4294_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na823_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y48     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4295_5 ( .OUT(na4295_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na843_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y51     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4296_5 ( .OUT(na4296_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na864_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y52     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4297_5 ( .OUT(na4297_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na864_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y53     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4298_5 ( .OUT(na4298_2), .IN1(1'b0), .IN2(na878_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x14y48     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4299_5 ( .OUT(na4299_2), .IN1(1'b0), .IN2(na878_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y49     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4300_5 ( .OUT(na4300_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na879_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y62     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4301_5 ( .OUT(na4301_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na880_2), .IN8(1'b0) );
// C_////Bridge      x44y51     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4302_5 ( .OUT(na4302_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na881_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y58     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4303_5 ( .OUT(na4303_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na884_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y51     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4304_5 ( .OUT(na4304_2), .IN1(1'b0), .IN2(1'b0), .IN3(na892_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4305_5 ( .OUT(na4305_2), .IN1(1'b0), .IN2(1'b0), .IN3(na892_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y58     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4306_5 ( .OUT(na4306_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na894_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y58     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4307_5 ( .OUT(na4307_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na894_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y50     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4308_5 ( .OUT(na4308_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na896_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y48     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4309_5 ( .OUT(na4309_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na896_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y44     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4310_5 ( .OUT(na4310_2), .IN1(1'b0), .IN2(na900_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y44     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4311_5 ( .OUT(na4311_2), .IN1(1'b0), .IN2(na900_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y39     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4312_5 ( .OUT(na4312_2), .IN1(1'b0), .IN2(na902_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y41     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4313_5 ( .OUT(na4313_2), .IN1(1'b0), .IN2(na902_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y45     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4314_5 ( .OUT(na4314_2), .IN1(1'b0), .IN2(na904_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y41     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4315_5 ( .OUT(na4315_2), .IN1(1'b0), .IN2(na904_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y43     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4316_5 ( .OUT(na4316_2), .IN1(1'b0), .IN2(na906_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y51     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4317_5 ( .OUT(na4317_2), .IN1(1'b0), .IN2(na906_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y46     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4318_5 ( .OUT(na4318_2), .IN1(na908_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y50     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4319_5 ( .OUT(na4319_2), .IN1(na908_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y42     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4320_5 ( .OUT(na4320_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na910_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y40     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4321_5 ( .OUT(na4321_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na910_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y46     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4322_5 ( .OUT(na4322_2), .IN1(1'b0), .IN2(na914_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y50     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4323_5 ( .OUT(na4323_2), .IN1(1'b0), .IN2(na914_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y42     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4324_5 ( .OUT(na4324_2), .IN1(1'b0), .IN2(1'b0), .IN3(na918_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y40     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4325_5 ( .OUT(na4325_2), .IN1(1'b0), .IN2(1'b0), .IN3(na918_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y43     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4326_5 ( .OUT(na4326_2), .IN1(1'b0), .IN2(na920_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y43     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4327_5 ( .OUT(na4327_2), .IN1(1'b0), .IN2(na920_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y40     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4328_5 ( .OUT(na4328_2), .IN1(1'b0), .IN2(1'b0), .IN3(na922_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y42     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4329_5 ( .OUT(na4329_2), .IN1(1'b0), .IN2(1'b0), .IN3(na922_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4330_5 ( .OUT(na4330_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na926_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y71     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4331_5 ( .OUT(na4331_2), .IN1(1'b0), .IN2(1'b0), .IN3(na928_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4332_5 ( .OUT(na4332_2), .IN1(1'b0), .IN2(1'b0), .IN3(na928_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y86     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4333_5 ( .OUT(na4333_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na986_1) );
// C_////Bridge      x41y84     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4334_5 ( .OUT(na4334_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na993_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4335_5 ( .OUT(na4335_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1010_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y75     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4336_5 ( .OUT(na4336_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1016_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y93     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4337_5 ( .OUT(na4337_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1038_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4338_5 ( .OUT(na4338_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1038_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y88     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4339_5 ( .OUT(na4339_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1043_1), .IN8(1'b0) );
// C_////Bridge      x48y88     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4340_5 ( .OUT(na4340_2), .IN1(1'b0), .IN2(na1044_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y71     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4341_5 ( .OUT(na4341_2), .IN1(1'b0), .IN2(na1052_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y73     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4342_5 ( .OUT(na4342_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1058_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y73     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4343_5 ( .OUT(na4343_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1058_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4344_5 ( .OUT(na4344_2), .IN1(na1062_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y72     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4345_5 ( .OUT(na4345_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1062_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y76     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4346_5 ( .OUT(na4346_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1064_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y78     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4347_5 ( .OUT(na4347_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1064_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4348_5 ( .OUT(na4348_2), .IN1(na1066_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y74     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4349_5 ( .OUT(na4349_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1066_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4350_5 ( .OUT(na4350_2), .IN1(na1068_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4351_5 ( .OUT(na4351_2), .IN1(na1068_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y74     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4352_5 ( .OUT(na4352_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1068_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4353_5 ( .OUT(na4353_2), .IN1(na1070_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y71     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4354_5 ( .OUT(na4354_2), .IN1(na1070_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y77     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4355_5 ( .OUT(na4355_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1072_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y75     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4356_5 ( .OUT(na4356_2), .IN1(na1072_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y75     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4357_5 ( .OUT(na4357_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1076_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y73     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4358_5 ( .OUT(na4358_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1076_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y76     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4359_5 ( .OUT(na4359_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1078_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y72     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4360_5 ( .OUT(na4360_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1078_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y69     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4361_5 ( .OUT(na4361_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1080_1) );
// C_////Bridge      x53y69     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4362_5 ( .OUT(na4362_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1080_2) );
// C_////Bridge      x55y76     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4363_5 ( .OUT(na4363_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1082_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4364_5 ( .OUT(na4364_2), .IN1(na1082_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4365_5 ( .OUT(na4365_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1090_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y74     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4366_5 ( .OUT(na4366_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1149_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4367_5 ( .OUT(na4367_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1149_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y85     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4368_5 ( .OUT(na4368_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1167_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y64     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4369_5 ( .OUT(na4369_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1179_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y89     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4370_5 ( .OUT(na4370_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1193_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y89     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4371_5 ( .OUT(na4371_2), .IN1(1'b0), .IN2(na1196_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y82     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4372_5 ( .OUT(na4372_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1198_1), .IN8(1'b0) );
// C_////Bridge      x51y78     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4373_5 ( .OUT(na4373_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1200_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y58     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4374_5 ( .OUT(na4374_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1200_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y62     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4375_5 ( .OUT(na4375_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1202_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y56     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4376_5 ( .OUT(na4376_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1202_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y60     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4377_5 ( .OUT(na4377_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1204_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y62     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4378_5 ( .OUT(na4378_2), .IN1(1'b0), .IN2(na1204_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y60     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4379_5 ( .OUT(na4379_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1208_1) );
// C_////Bridge      x35y58     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4380_5 ( .OUT(na4380_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1208_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y66     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4381_5 ( .OUT(na4381_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1210_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x30y66     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4382_5 ( .OUT(na4382_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1210_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4383_5 ( .OUT(na4383_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1212_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4384_5 ( .OUT(na4384_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1212_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y61     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4385_5 ( .OUT(na4385_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1214_1) );
// C_////Bridge      x36y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4386_5 ( .OUT(na4386_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1214_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4387_5 ( .OUT(na4387_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1216_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y57     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4388_5 ( .OUT(na4388_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1216_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y62     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4389_5 ( .OUT(na4389_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1222_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y62     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4390_5 ( .OUT(na4390_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1222_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4391_5 ( .OUT(na4391_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1224_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y58     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4392_5 ( .OUT(na4392_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1226_1), .IN8(1'b0) );
// C_////Bridge      x34y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4393_5 ( .OUT(na4393_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1226_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y57     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4394_5 ( .OUT(na4394_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1228_1) );
// C_////Bridge      x38y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4395_5 ( .OUT(na4395_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1228_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y54     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4396_5 ( .OUT(na4396_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1230_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y54     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4397_5 ( .OUT(na4397_2), .IN1(na1230_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y84     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4398_5 ( .OUT(na4398_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1260_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y73     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4399_5 ( .OUT(na4399_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1296_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4400_5 ( .OUT(na4400_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1296_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y74     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4401_5 ( .OUT(na4401_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1296_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y88     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4402_5 ( .OUT(na4402_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1306_1) );
// C_////Bridge      x31y81     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4403_5 ( .OUT(na4403_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1313_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y87     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4404_5 ( .OUT(na4404_2), .IN1(1'b0), .IN2(na1321_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y89     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4405_5 ( .OUT(na4405_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1324_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y87     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4406_5 ( .OUT(na4406_2), .IN1(1'b0), .IN2(na1325_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y85     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4407_5 ( .OUT(na4407_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1326_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4408_5 ( .OUT(na4408_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1330_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y69     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4409_5 ( .OUT(na4409_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1330_2) );
// C_////Bridge      x31y85     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4410_5 ( .OUT(na4410_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1331_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x43y89     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4411_5 ( .OUT(na4411_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1347_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y92     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4412_5 ( .OUT(na4412_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1349_2), .IN8(1'b0) );
// C_////Bridge      x11y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4413_5 ( .OUT(na4413_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1351_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y41     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4414_5 ( .OUT(na4414_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1353_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y68     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4415_5 ( .OUT(na4415_2), .IN1(na1366_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y56     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4416_5 ( .OUT(na4416_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1375_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y85     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4417_5 ( .OUT(na4417_2), .IN1(1'b0), .IN2(na1377_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y54     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4418_5 ( .OUT(na4418_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1386_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y63     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4419_5 ( .OUT(na4419_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1387_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y73     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4420_5 ( .OUT(na4420_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1438_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x69y80     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4421_5 ( .OUT(na4421_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1439_1), .IN8(1'b0) );
// C_////Bridge      x57y83     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4422_5 ( .OUT(na4422_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1440_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y65     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4423_5 ( .OUT(na4423_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1443_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y64     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4424_5 ( .OUT(na4424_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1443_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x69y70     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4425_5 ( .OUT(na4425_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1444_1), .IN8(1'b0) );
// C_////Bridge      x71y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4426_5 ( .OUT(na4426_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1446_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4427_5 ( .OUT(na4427_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1447_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y73     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4428_5 ( .OUT(na4428_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1451_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y57     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4429_5 ( .OUT(na4429_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1460_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y67     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4430_5 ( .OUT(na4430_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1461_1) );
// C_////Bridge      x55y74     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4431_5 ( .OUT(na4431_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1462_2), .IN8(1'b0) );
// C_////Bridge      x54y50     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4432_5 ( .OUT(na4432_2), .IN1(na1465_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y53     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4433_5 ( .OUT(na4433_2), .IN1(1'b0), .IN2(na1466_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y58     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4434_5 ( .OUT(na4434_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1467_2), .IN8(1'b0) );
// C_////Bridge      x57y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4435_5 ( .OUT(na4435_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1468_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y48     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4436_5 ( .OUT(na4436_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1469_1), .IN8(1'b0) );
// C_////Bridge      x50y62     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4437_5 ( .OUT(na4437_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1473_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y55     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4438_5 ( .OUT(na4438_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1482_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y66     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4439_5 ( .OUT(na4439_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1483_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x18y72     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4440_5 ( .OUT(na4440_2), .IN1(na1484_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x15y48     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4441_5 ( .OUT(na4441_2), .IN1(1'b0), .IN2(na1487_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y52     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4442_5 ( .OUT(na4442_2), .IN1(1'b0), .IN2(na1487_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y64     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4443_5 ( .OUT(na4443_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1488_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y47     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4444_5 ( .OUT(na4444_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1489_2) );
// C_////Bridge      x20y50     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4445_5 ( .OUT(na4445_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1490_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y54     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4446_5 ( .OUT(na4446_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1491_1), .IN8(1'b0) );
// C_////Bridge      x42y87     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4447_5 ( .OUT(na4447_2), .IN1(1'b0), .IN2(na1504_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y89     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4448_5 ( .OUT(na4448_2), .IN1(1'b0), .IN2(na1505_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x30y91     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4449_5 ( .OUT(na4449_2), .IN1(1'b0), .IN2(na1506_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y90     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4450_5 ( .OUT(na4450_2), .IN1(na1510_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y87     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4451_5 ( .OUT(na4451_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1512_1) );
// C_////Bridge      x34y81     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4452_5 ( .OUT(na4452_2), .IN1(1'b0), .IN2(na1513_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y85     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4453_5 ( .OUT(na4453_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1526_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y92     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4454_5 ( .OUT(na4454_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1527_2), .IN8(1'b0) );
// C_////Bridge      x50y91     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4455_5 ( .OUT(na4455_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1528_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4456_5 ( .OUT(na4456_2), .IN1(na1532_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y92     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4457_5 ( .OUT(na4457_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1533_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y86     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4458_5 ( .OUT(na4458_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1534_2), .IN8(1'b0) );
// C_////Bridge      x64y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4459_5 ( .OUT(na4459_2), .IN1(na1535_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y61     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4460_5 ( .OUT(na4460_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1539_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y61     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4461_5 ( .OUT(na4461_2), .IN1(1'b0), .IN2(na1541_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y60     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4462_5 ( .OUT(na4462_2), .IN1(1'b0), .IN2(na1541_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y40     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4463_5 ( .OUT(na4463_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1542_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y37     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4464_5 ( .OUT(na4464_2), .IN1(1'b0), .IN2(na1542_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4465_5 ( .OUT(na4465_2), .IN1(1'b0), .IN2(na1543_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4466_5 ( .OUT(na4466_2), .IN1(1'b0), .IN2(na1543_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y47     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4467_5 ( .OUT(na4467_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1544_2) );
// C_////Bridge      x41y45     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4468_5 ( .OUT(na4468_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1545_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x15y56     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4469_5 ( .OUT(na4469_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1567_2), .IN8(1'b0) );
// C_////Bridge      x15y63     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4470_5 ( .OUT(na4470_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1610_1) );
// C_////Bridge      x13y63     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4471_5 ( .OUT(na4471_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1610_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x12y63     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4472_5 ( .OUT(na4472_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1610_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y67     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4473_5 ( .OUT(na4473_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1613_1), .IN8(1'b0) );
// C_////Bridge      x16y65     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4474_5 ( .OUT(na4474_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1614_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y65     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4475_5 ( .OUT(na4475_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1771_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y66     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4476_5 ( .OUT(na4476_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1773_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y65     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4477_5 ( .OUT(na4477_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1773_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y48     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4478_5 ( .OUT(na4478_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1811_1), .IN8(1'b0) );
// C_////Bridge      x30y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4479_5 ( .OUT(na4479_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1811_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y58     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4480_5 ( .OUT(na4480_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1864_1), .IN8(1'b0) );
// C_////Bridge      x64y51     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4481_5 ( .OUT(na4481_2), .IN1(na1887_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y53     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4482_5 ( .OUT(na4482_2), .IN1(na1887_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x69y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4483_5 ( .OUT(na4483_2), .IN1(1'b0), .IN2(na1986_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y66     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4484_5 ( .OUT(na4484_2), .IN1(1'b0), .IN2(na1986_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4485_5 ( .OUT(na4485_2), .IN1(1'b0), .IN2(na1986_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x72y72     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4486_5 ( .OUT(na4486_2), .IN1(1'b0), .IN2(na1986_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y71     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4487_5 ( .OUT(na4487_2), .IN1(1'b0), .IN2(na1989_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y69     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4488_5 ( .OUT(na4488_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1990_1) );
// C_////Bridge      x65y67     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4489_5 ( .OUT(na4489_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1990_2) );
// C_////Bridge      x67y67     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4490_5 ( .OUT(na4490_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1991_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y67     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4491_5 ( .OUT(na4491_2), .IN1(1'b0), .IN2(na1993_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y74     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4492_5 ( .OUT(na4492_2), .IN1(1'b0), .IN2(na1993_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y61     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4493_5 ( .OUT(na4493_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1993_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y49     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4494_5 ( .OUT(na4494_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na1999_1), .IN8(1'b0) );
// C_////Bridge      x49y49     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4495_5 ( .OUT(na4495_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2000_2) );
// C_////Bridge      x47y51     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4496_5 ( .OUT(na4496_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2002_1), .IN8(1'b0) );
// C_////Bridge      x54y56     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4497_5 ( .OUT(na4497_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2013_2), .IN8(1'b0) );
// C_////Bridge      x56y57     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4498_5 ( .OUT(na4498_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2015_1) );
// C_////Bridge      x52y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4499_5 ( .OUT(na4499_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2017_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y51     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4500_5 ( .OUT(na4500_2), .IN1(na2122_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y55     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4501_5 ( .OUT(na4501_2), .IN1(na2122_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y63     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4502_5 ( .OUT(na4502_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2124_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x66y52     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4503_5 ( .OUT(na4503_2), .IN1(na2222_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y56     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4504_5 ( .OUT(na4504_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2223_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x65y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4505_5 ( .OUT(na4505_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2226_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y61     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4506_5 ( .OUT(na4506_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2228_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y63     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4507_5 ( .OUT(na4507_2), .IN1(1'b0), .IN2(na2228_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y60     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4508_5 ( .OUT(na4508_2), .IN1(1'b0), .IN2(na2228_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y58     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4509_5 ( .OUT(na4509_2), .IN1(na2229_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y64     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4510_5 ( .OUT(na4510_2), .IN1(na2229_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y62     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4511_5 ( .OUT(na4511_2), .IN1(na2229_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y57     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4512_5 ( .OUT(na4512_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2230_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y46     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4513_5 ( .OUT(na4513_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2236_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y52     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4514_5 ( .OUT(na4514_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2237_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y50     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4515_5 ( .OUT(na4515_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2239_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y56     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4516_5 ( .OUT(na4516_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2250_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y54     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4517_5 ( .OUT(na4517_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2252_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y51     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4518_5 ( .OUT(na4518_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2254_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x70y67     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4519_5 ( .OUT(na4519_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2350_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4520_5 ( .OUT(na4520_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2473_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y65     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4521_5 ( .OUT(na4521_2), .IN1(1'b0), .IN2(na2474_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y53     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4522_5 ( .OUT(na4522_2), .IN1(1'b0), .IN2(na2474_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y55     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4523_5 ( .OUT(na4523_2), .IN1(1'b0), .IN2(na2474_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y55     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4524_5 ( .OUT(na4524_2), .IN1(1'b0), .IN2(na2477_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x18y56     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4525_5 ( .OUT(na4525_2), .IN1(1'b0), .IN2(na2477_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y51     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4526_5 ( .OUT(na4526_2), .IN1(1'b0), .IN2(na2478_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y56     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4527_5 ( .OUT(na4527_2), .IN1(1'b0), .IN2(na2478_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y61     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4528_5 ( .OUT(na4528_2), .IN1(1'b0), .IN2(na2478_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y55     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4529_5 ( .OUT(na4529_2), .IN1(1'b0), .IN2(na2478_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y53     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4530_5 ( .OUT(na4530_2), .IN1(1'b0), .IN2(na2478_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y48     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4531_5 ( .OUT(na4531_2), .IN1(na2479_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x20y56     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4532_5 ( .OUT(na4532_2), .IN1(na2479_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x19y50     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4533_5 ( .OUT(na4533_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2481_1), .IN8(1'b0) );
// C_////Bridge      x23y45     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4534_5 ( .OUT(na4534_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2481_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y52     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4535_5 ( .OUT(na4535_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2481_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y38     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4536_5 ( .OUT(na4536_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2487_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y34     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4537_5 ( .OUT(na4537_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2488_1), .IN8(1'b0) );
// C_////Bridge      x22y36     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4538_5 ( .OUT(na4538_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2490_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y44     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4539_5 ( .OUT(na4539_2), .IN1(na2501_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y45     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4540_5 ( .OUT(na4540_2), .IN1(1'b0), .IN2(na2503_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x17y42     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4541_5 ( .OUT(na4541_2), .IN1(na2505_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y60     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4542_5 ( .OUT(na4542_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2529_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y45     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4543_5 ( .OUT(na4543_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2599_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y84     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4544_5 ( .OUT(na4544_2), .IN1(1'b0), .IN2(na2706_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y91     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4545_5 ( .OUT(na4545_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2707_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y86     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4546_5 ( .OUT(na4546_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2707_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y83     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4547_5 ( .OUT(na4547_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2707_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y91     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4548_5 ( .OUT(na4548_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2707_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y80     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4549_5 ( .OUT(na4549_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2712_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y84     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4550_5 ( .OUT(na4550_2), .IN1(na2712_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4551_5 ( .OUT(na4551_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2713_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4552_5 ( .OUT(na4552_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2713_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y82     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4553_5 ( .OUT(na4553_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2713_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4554_5 ( .OUT(na4554_2), .IN1(na2714_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y67     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4555_5 ( .OUT(na4555_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2720_1) );
// C_////Bridge      x37y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4556_5 ( .OUT(na4556_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2721_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y69     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4557_5 ( .OUT(na4557_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2722_2) );
// C_////Bridge      x57y87     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4558_5 ( .OUT(na4558_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na2730_2) );
// C_////Bridge      x33y67     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4559_5 ( .OUT(na4559_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2741_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y69     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4560_5 ( .OUT(na4560_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2743_2), .IN8(1'b0) );
// C_////Bridge      x27y73     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4561_5 ( .OUT(na4561_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2745_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y76     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4562_5 ( .OUT(na4562_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na2846_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4563_5 ( .OUT(na4563_2), .IN1(na2957_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y84     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4564_5 ( .OUT(na4564_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2958_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x68y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4565_5 ( .OUT(na4565_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2958_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y86     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4566_5 ( .OUT(na4566_2), .IN1(1'b0), .IN2(1'b0), .IN3(na2958_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y84     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4567_5 ( .OUT(na4567_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na2961_1), .IN8(1'b0) );
// C_////Bridge      x60y84     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4568_5 ( .OUT(na4568_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2962_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y84     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4569_5 ( .OUT(na4569_2), .IN1(na2962_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y81     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4570_5 ( .OUT(na4570_2), .IN1(na2962_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y86     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4571_5 ( .OUT(na4571_2), .IN1(na2962_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4572_5 ( .OUT(na4572_2), .IN1(na2963_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y83     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4573_5 ( .OUT(na4573_2), .IN1(1'b0), .IN2(na2965_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x16y62     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4574_5 ( .OUT(na4574_2), .IN1(1'b0), .IN2(na2973_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y64     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4575_5 ( .OUT(na4575_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2973_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y60     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4576_5 ( .OUT(na4576_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na2974_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y73     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4577_5 ( .OUT(na4577_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na2981_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y66     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4578_5 ( .OUT(na4578_2), .IN1(na2988_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4579_5 ( .OUT(na4579_2), .IN1(1'b0), .IN2(na2990_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y76     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4580_5 ( .OUT(na4580_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3104_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y76     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4581_5 ( .OUT(na4581_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3230_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x18y63     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4582_5 ( .OUT(na4582_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na3258_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y64     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4583_5 ( .OUT(na4583_2), .IN1(na3278_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y64     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4584_5 ( .OUT(na4584_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3282_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x71y49     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4585_5 ( .OUT(na4585_2), .IN1(1'b0), .IN2(na3283_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y42     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4586_5 ( .OUT(na4586_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3288_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y47     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4587_5 ( .OUT(na4587_2), .IN1(na3303_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y61     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4588_5 ( .OUT(na4588_2), .IN1(1'b0), .IN2(na3313_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y88     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4589_5 ( .OUT(na4589_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3329_2) );
// C_////Bridge      x69y81     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4590_5 ( .OUT(na4590_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3348_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y74     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4591_5 ( .OUT(na4591_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3416_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y70     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4592_5 ( .OUT(na4592_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3417_1), .IN8(1'b0) );
// C_////Bridge      x58y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4593_5 ( .OUT(na4593_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3423_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y74     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4594_5 ( .OUT(na4594_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3424_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y52     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4595_5 ( .OUT(na4595_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3426_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y52     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4596_5 ( .OUT(na4596_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3427_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y58     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4597_5 ( .OUT(na4597_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3429_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y54     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4598_5 ( .OUT(na4598_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3430_1), .IN8(1'b0) );
// C_////Bridge      x35y60     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4599_5 ( .OUT(na4599_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3439_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y58     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4600_5 ( .OUT(na4600_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3442_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y56     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4601_5 ( .OUT(na4601_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3443_2), .IN8(1'b0) );
// C_////Bridge      x33y56     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4602_5 ( .OUT(na4602_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3444_1), .IN8(1'b0) );
// C_////Bridge      x66y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4603_5 ( .OUT(na4603_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3451_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y54     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4604_5 ( .OUT(na4604_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3472_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y39     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4605_5 ( .OUT(na4605_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3525_2) );
// C_////Bridge      x42y41     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4606_5 ( .OUT(na4606_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3526_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y41     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4607_5 ( .OUT(na4607_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3529_2) );
// C_////Bridge      x44y41     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4608_5 ( .OUT(na4608_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3530_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y73     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4609_5 ( .OUT(na4609_2), .IN1(na3578_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y73     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4610_5 ( .OUT(na4610_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3580_1), .IN8(1'b0) );
// C_////Bridge      x18y51     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4611_5 ( .OUT(na4611_2), .IN1(na3590_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y88     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4612_5 ( .OUT(na4612_2), .IN1(1'b0), .IN2(na3701_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y85     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4613_5 ( .OUT(na4613_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3708_2), .IN8(1'b0) );
// C_////Bridge      x64y45     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4614_5 ( .OUT(na4614_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3711_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x64y43     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4615_5 ( .OUT(na4615_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3712_1) );
// C_////Bridge      x58y41     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4616_5 ( .OUT(na4616_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3715_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y41     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4617_5 ( .OUT(na4617_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3716_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y34     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4618_5 ( .OUT(na4618_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3719_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y34     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4619_5 ( .OUT(na4619_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3720_1) );
// C_////Bridge      x65y36     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4620_5 ( .OUT(na4620_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3721_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x63y40     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4621_5 ( .OUT(na4621_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3722_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y36     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4622_5 ( .OUT(na4622_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na3723_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y36     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4623_5 ( .OUT(na4623_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na3724_1) );
// C_////Bridge      x67y36     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4624_5 ( .OUT(na4624_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3725_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x67y34     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4625_5 ( .OUT(na4625_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3726_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y88     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4626_5 ( .OUT(na4626_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na3815_1), .IN8(1'b0) );
// C_////Bridge      x64y92     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4627_5 ( .OUT(na4627_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3828_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y60     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4628_5 ( .OUT(na4628_2), .IN1(1'b0), .IN2(1'b0), .IN3(na3898_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y87     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4629_5 ( .OUT(na4629_2), .IN1(na3931_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y92     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4630_5 ( .OUT(na4630_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na3931_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y79     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4631_5 ( .OUT(na4631_2), .IN1(1'b0), .IN2(na3943_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a4632_5 ( .OUT(na4632_2), .IN1(1'b0), .IN2(na3943_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
endmodule
