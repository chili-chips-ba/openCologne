//  (c) Cologne Chip AG
//  FPGA Verilog netlist writer     Version: Version 4.2 (1 July 2024)
//  Compile Time: 2024-07-19 13:57:40
//  Program Run:  2024-08-04 23:01:36
//  Program Call: /home/user/FPGA/Boards/GateMate/cc-toolchain-linux//bin/p_r/p_r -i net/fm_synth.v -o fm -ccf fm.ccf -cCP 
//  File Type:    Verilog

// Gatecount:   1325
module fm (btn , clk_10mhz ,
       ant_433mhz , led , wifi_gpio0 
       ) ;

input  btn;
input  clk_10mhz;

output ant_433mhz;
output led;
output wifi_gpio0;



wire btn;
wire led;
wire na4_1;
wire na5_2;
wire na6_1;
wire na7_2;
wire na8_1;
wire na9_1;
wire na10_1;
wire na11_1;
wire na12_1;
wire na13_1;
wire na14_1;
wire na15_1;
wire na16_1;
wire na17_1;
wire na18_1;
wire na19_2;
wire na20_2;
wire na21_2;
wire na22_1;
wire na23_2;
wire na24_1;
wire na24_2;
wire na25_1;
wire na26_2;
wire na27_1;
wire na28_1;
wire na29_2;
wire na30_1;
wire na31_2;
wire na32_1;
wire na32_2;
wire na35_1;
wire na35_1_i;
wire na36_1;
wire na36_1_i;
wire na37_1;
wire na37_1_i;
wire na38_1;
wire na38_1_i;
wire na39_1;
wire na39_1_i;
wire na40_1;
wire na40_1_i;
wire na41_1;
wire na41_1_i;
wire na42_1;
wire na42_1_i;
wire na43_1;
wire na43_1_i;
wire na44_1;
wire na44_1_i;
wire na45_1;
wire na45_1_i;
wire na46_1;
wire na46_1_i;
wire na47_1;
wire na47_1_i;
wire na48_1;
wire na48_1_i;
wire na49_1;
wire na49_1_i;
wire na50_1;
wire na50_2;
wire na51_1;
wire na52_2;
wire na53_1;
wire na54_1;
wire na55_1;
wire na56_1;
wire na57_1;
wire na58_2;
wire na60_1;
wire na61_1;
wire na62_1;
wire na63_1;
wire na64_2;
wire na65_1;
wire na66_1;
wire na67_1;
wire na68_1;
wire na69_1;
wire na70_1;
wire na72_2;
wire na72_2_i;
wire na73_1;
wire na73_1_i;
wire na74_1;
wire na74_1_i;
wire na75_1;
wire na75_1_i;
wire na76_1;
wire na76_1_i;
wire na77_1;
wire na77_1_i;
wire na78_1;
wire na78_1_i;
wire na79_1;
wire na79_1_i;
wire na80_1;
wire na80_1_i;
wire na81_1;
wire na81_1_i;
wire na82_1;
wire na82_1_i;
wire na83_1;
wire na83_1_i;
wire na84_2;
wire na85_1;
wire na85_1_i;
wire na86_1;
wire na86_1_i;
wire na87_1;
wire na87_1_i;
wire na88_1;
wire na88_1_i;
wire na89_1;
wire na89_1_i;
wire na90_1;
wire na90_1_i;
wire na91_1;
wire na91_1_i;
wire na91_2;
wire na91_2_i;
wire na93_1;
wire na93_1_i;
wire na94_2;
wire na94_2_i;
wire na95_1;
wire na97_1;
wire na97_1_i;
wire na98_1;
wire na98_1_i;
wire na98_2;
wire na98_2_i;
wire na99_1;
wire na99_1_i;
wire na99_2;
wire na99_2_i;
wire na103_1;
wire na106_2;
wire na106_2_i;
wire na107_1;
wire na107_1_i;
wire na108_2;
wire na108_2_i;
wire na109_1;
wire na109_1_i;
wire na109_2;
wire na109_2_i;
wire na110_1;
wire na110_1_i;
wire na110_2;
wire na110_2_i;
wire na111_1;
wire na111_1_i;
wire na112_1;
wire na112_1_i;
wire na113_2;
wire na113_2_i;
wire na114_1;
wire na114_1_i;
wire na115_2;
wire na115_2_i;
wire na116_1;
wire na116_1_i;
wire na116_2;
wire na116_2_i;
wire na118_1;
wire na118_1_i;
wire na119_2;
wire na119_2_i;
wire na120_1;
wire na121_1;
wire na122_1;
wire na124_2;
wire na125_2;
wire na127_1;
wire na128_1;
wire na128_2;
wire na129_2;
wire na131_1;
wire na132_1;
wire na132_2;
wire na133_2;
wire na135_1;
wire na136_1;
wire na136_2;
wire na137_2;
wire na138_1;
wire na139_1;
wire na140_1;
wire na142_1;
wire na143_1;
wire na145_2;
wire na146_1;
wire na146_2;
wire na147_1;
wire na149_2;
wire na150_1;
wire na150_2;
wire na151_1;
wire na153_2;
wire na154_1;
wire na154_2;
wire na155_1;
wire na156_1;
wire na157_1;
wire na161_1;
wire na161_2;
wire na162_2;
wire na164_1;
wire na165_1;
wire na166_1;
wire na166_1_i;
wire na167_1;
wire na168_1;
wire na169_1;
wire na171_2;
wire na172_2;
wire na173_1;
wire na173_2;
wire na176_1;
wire na176_2;
wire na177_1;
wire na178_1;
wire na179_1;
wire na180_1;
wire na181_1;
wire na182_1;
wire na184_1;
wire na185_2;
wire na186_1;
wire na187_1;
wire na188_1;
wire na189_2;
wire na190_1;
wire na191_2;
wire na192_1;
wire na193_1;
wire na194_1;
wire na195_1;
wire na196_1;
wire na197_1;
wire na198_1;
wire na199_1;
wire na200_2;
wire na201_1;
wire na202_1;
wire na203_1;
wire na204_1;
wire na205_1;
wire na206_1;
wire na207_2;
wire na208_1;
wire na209_2;
wire na210_1;
wire na211_1;
wire na212_1;
wire na213_1;
wire na214_1;
wire na215_1;
wire na216_1;
wire na217_1;
wire na218_2;
wire na219_1;
wire na220_1;
wire na221_1;
wire na222_1;
wire na223_1;
wire na224_1;
wire na225_2;
wire na226_1;
wire na227_2;
wire na228_1;
wire na229_1;
wire na230_1;
wire na231_1;
wire na232_1;
wire na233_1;
wire na234_2;
wire na235_1;
wire na236_2;
wire na237_1;
wire na238_1;
wire na239_1;
wire na240_1;
wire na241_2;
wire na242_1;
wire na243_1;
wire na244_1;
wire na245_2;
wire na246_1;
wire na247_1;
wire na248_2;
wire na249_1;
wire na250_1;
wire na251_1;
wire na251_2;
wire na252_1;
wire na252_2;
wire na254_1;
wire na254_2;
wire na256_1;
wire na256_2;
wire na258_1;
wire na258_2;
wire na259_2;
wire na260_1;
wire na261_1;
wire na262_1;
wire na265_1;
wire na267_1;
wire na269_1;
wire na272_1;
wire na274_1;
wire na275_1;
wire na275_2;
wire na277_1;
wire na279_1;
wire na282_1;
wire na284_1;
wire na285_2;
wire na288_1;
wire na290_1;
wire na290_2;
wire na292_1;
wire na292_2;
wire na293_1;
wire na295_1;
wire na296_1;
wire na297_1;
wire na298_1;
wire na299_1;
wire na300_1;
wire na301_1;
wire na302_2;
wire na303_1;
wire na304_2;
wire na305_1;
wire na307_1;
wire na307_2;
wire na309_1;
wire na309_2;
wire na311_1;
wire na311_2;
wire na312_2;
wire na314_1;
wire na318_1;
wire na319_1;
wire na321_1;
wire na322_2;
wire na323_1;
wire na324_1;
wire na325_1;
wire na326_1;
wire na327_2;
wire na328_1;
wire na329_1;
wire na330_2;
wire na331_1;
wire na333_1;
wire na333_2;
wire na335_1;
wire na335_2;
wire na337_1;
wire na337_2;
wire na338_2;
wire na340_1;
wire na344_1;
wire na345_1;
wire na411_4;
wire na413_4;
wire na414_2;
wire na414_4;
wire na415_1;
wire na415_4;
wire na416_4;
wire na418_4;
wire na420_4;
wire na422_4;
wire na424_4;
wire na425_1;
wire na425_4;
wire na426_1;
wire na426_1_i;
wire na426_2;
wire na428_1;
wire na428_4;
wire na429_1;
wire na429_1_i;
wire na429_2;
wire na429_4;
wire na431_1;
wire na431_1_i;
wire na431_2;
wire na433_1;
wire na433_4;
wire na434_1;
wire na434_2;
wire na434_4;
wire na436_1;
wire na436_2;
wire na437_1;
wire na437_4;
wire na439_1;
wire na439_2;
wire na439_4;
wire na441_1;
wire na441_2;
wire na441_4;
wire na443_1;
wire na444_1;
wire na444_2;
wire na444_4;
wire na446_1;
wire na446_2;
wire na446_4;
wire na448_1;
wire na448_2;
wire na448_4;
wire na450_1;
wire na450_2;
wire na450_4;
wire na452_1;
wire na452_2;
wire na452_4;
wire na453_1;
wire na453_4;
wire na455_1;
wire na455_2;
wire na455_4;
wire na457_1;
wire na457_2;
wire na457_4;
wire na459_1;
wire na460_1;
wire na460_2;
wire na460_4;
wire na462_1;
wire na462_2;
wire na462_4;
wire na464_1;
wire na464_2;
wire na464_4;
wire na466_1;
wire na466_2;
wire na466_4;
wire na468_1;
wire na468_2;
wire na468_4;
wire na469_1;
wire na469_4;
wire na471_1;
wire na471_1_i;
wire na471_2;
wire na471_4;
wire na473_1;
wire na473_1_i;
wire na473_2;
wire na473_4;
wire na475_1;
wire na475_1_i;
wire na475_2;
wire na475_4;
wire na477_1;
wire na477_1_i;
wire na477_2;
wire na477_4;
wire na479_1;
wire na479_1_i;
wire na479_2;
wire na479_4;
wire na480_1;
wire na480_1_i;
wire na480_2;
wire na480_4;
wire na482_1;
wire na482_1_i;
wire na482_2;
wire na482_4;
wire na484_1;
wire na484_1_i;
wire na484_2;
wire na484_4;
wire na486_1;
wire na486_1_i;
wire na486_2;
wire na489_1;
wire na489_1_i;
wire na489_2;
wire na489_4;
wire na491_1;
wire na491_1_i;
wire na491_2;
wire na491_4;
wire na493_1;
wire na493_1_i;
wire na493_2;
wire na493_4;
wire na495_1;
wire na495_1_i;
wire na495_2;
wire na495_4;
wire na496_1;
wire na496_4;
wire na498_1;
wire na498_1_i;
wire na498_2;
wire na498_4;
wire na500_1;
wire na500_1_i;
wire na500_2;
wire na500_4;
wire na502_1;
wire na502_1_i;
wire na503_1;
wire na503_1_i;
wire na503_2;
wire na503_4;
wire na505_1;
wire na505_1_i;
wire na505_2;
wire na505_4;
wire na507_1;
wire na507_1_i;
wire na507_2;
wire na507_4;
wire na509_1;
wire na509_1_i;
wire na509_2;
wire na509_4;
wire na511_1;
wire na511_1_i;
wire na511_2;
wire na511_4;
wire na512_1;
wire na512_1_i;
wire na512_2;
wire na512_4;
wire na513_1;
wire na513_1_i;
wire na513_2;
wire na513_4;
wire na515_1;
wire na515_1_i;
wire na515_2;
wire na515_4;
wire na517_1;
wire na517_1_i;
wire na517_2;
wire na517_4;
wire na519_1;
wire na519_1_i;
wire na519_2;
wire na519_4;
wire na521_1;
wire na521_1_i;
wire na521_2;
wire na521_4;
wire na524_1;
wire na524_1_i;
wire na524_2;
wire na524_4;
wire na526_1;
wire na526_1_i;
wire na526_2;
wire na526_4;
wire na528_1;
wire na528_1_i;
wire na528_2;
wire na528_4;
wire na530_1;
wire na530_1_i;
wire na530_2;
wire na532_1;
wire na532_1_i;
wire na532_2;
wire na532_4;
wire na534_1;
wire na534_1_i;
wire na534_2;
wire na534_4;
wire na536_1;
wire na536_1_i;
wire na536_2;
wire na536_4;
wire na538_1;
wire na538_1_i;
wire na538_2;
wire na538_4;
wire na540_1;
wire na540_4;
wire na541_1;
wire na541_2;
wire na541_4;
wire na543_1;
wire na543_2;
wire na543_4;
wire na545_1;
wire na546_1;
wire na546_4;
wire na547_1;
wire na547_2;
wire na547_4;
wire na549_1;
wire na549_2;
wire na549_4;
wire na551_1;
wire na552_1;
wire na552_4;
wire na553_1;
wire na553_2;
wire na553_4;
wire na555_1;
wire na555_2;
wire na555_4;
wire na557_1;
wire na557_2;
wire na559_1;
wire na559_2;
wire na559_4;
wire na560_1;
wire na560_2;
wire na560_4;
wire na562_1;
wire na562_2;
wire na562_4;
wire na564_1;
wire na564_2;
wire na567_1;
wire na567_2;
wire na567_4;
wire na569_1;
wire na569_2;
wire na569_4;
wire na571_1;
wire na571_2;
wire na571_4;
wire na573_1;
wire na573_2;
wire na573_4;
wire na575_1;
wire na575_4;
wire na576_1;
wire na576_2;
wire na576_4;
wire na578_1;
wire na578_2;
wire na578_4;
wire na580_1;
wire na580_4;
wire na581_1;
wire na581_4;
wire na582_1;
wire na582_4;
wire na583_1;
wire na583_1_i;
wire na583_2;
wire na583_4;
wire na585_1;
wire na585_1_i;
wire na585_2;
wire na587_1;
wire na587_4;
wire na589_1;
wire na590_1;
wire na590_2;
wire na590_4;
wire na592_1;
wire na592_2;
wire na592_4;
wire na594_1;
wire na594_2;
wire na594_4;
wire na596_1;
wire na596_2;
wire na596_4;
wire na598_1;
wire na598_2;
wire na598_4;
wire na599_1;
wire na599_4;
wire na601_1;
wire na601_2;
wire na601_4;
wire na603_1;
wire na603_2;
wire na603_4;
wire na605_1;
wire na605_2;
wire na605_4;
wire na607_1;
wire na607_2;
wire na607_4;
wire na609_1;
wire na609_2;
wire na610_1;
wire na610_4;
wire na611_1;
wire na611_1_i;
wire na611_2;
wire na611_4;
wire na613_1;
wire na613_1_i;
wire na613_2;
wire na615_1;
wire na615_4;
wire na616_1;
wire na616_2;
wire na616_4;
wire na618_1;
wire na618_2;
wire na618_4;
wire na620_1;
wire na620_4;
wire na621_1;
wire na621_4;
wire na624_1;
wire na624_2;
wire na634_2;
wire na634_2_i;
wire na635_1;
wire na635_1_i;
wire na636_1;
wire na636_1_i;
wire na638_1;
wire na638_1_i;
wire na640_2;
wire na640_2_i;
wire na642_1;
wire na642_1_i;
wire na644_2;
wire na644_2_i;
wire na646_1;
wire na646_1_i;
wire na648_2;
wire na648_2_i;
wire na650_1;
wire na650_1_i;
wire na652_2;
wire na652_2_i;
wire na654_1;
wire na654_1_i;
wire na656_2;
wire na656_2_i;
wire na658_1;
wire na658_1_i;
wire na660_2;
wire na660_2_i;
wire na662_1;
wire na662_1_i;
wire na663_2;
wire na663_2_i;
wire na696_1;
wire na696_1_i;
wire na696_2;
wire na696_2_i;
wire na698_1;
wire na698_1_i;
wire na700_2;
wire na700_2_i;
wire na702_1;
wire na702_1_i;
wire na704_2;
wire na704_2_i;
wire na706_1;
wire na706_1_i;
wire na708_2;
wire na708_2_i;
wire na720_1;
wire na720_1_i;
wire na721_1;
wire na721_1_i;
wire na721_2;
wire na721_2_i;
wire na722_2;
wire na722_2_i;
wire na723_1;
wire na723_1_i;
wire na723_2;
wire na723_2_i;
wire na724_1;
wire na724_1_i;
wire na725_1;
wire na725_1_i;
wire na725_2;
wire na725_2_i;
wire na726_2;
wire na726_2_i;
wire na727_1;
wire na727_1_i;
wire na727_2;
wire na727_2_i;
wire na728_1;
wire na728_1_i;
wire na729_1;
wire na729_1_i;
wire na729_2;
wire na729_2_i;
wire na730_1;
wire na730_1_i;
wire na731_1;
wire na731_1_i;
wire na731_2;
wire na731_2_i;
wire na732_2;
wire na732_2_i;
wire na733_1;
wire na733_1_i;
wire na733_2;
wire na733_2_i;
wire na734_1;
wire na734_1_i;
wire na734_2;
wire na734_2_i;
wire na735_1;
wire na735_1_i;
wire na744_2;
wire na744_2_i;
wire na745_1;
wire na745_1_i;
wire na745_2;
wire na745_2_i;
wire na748_1;
wire na748_1_i;
wire na750_2;
wire na750_2_i;
wire na752_1;
wire na752_1_i;
wire na754_1;
wire na754_1_i;
wire na756_2;
wire na756_2_i;
wire na758_2;
wire na758_2_i;
wire na760_2;
wire na760_2_i;
wire na762_1;
wire na762_1_i;
wire na764_2;
wire na764_2_i;
wire na766_1;
wire na766_1_i;
wire na768_1;
wire na768_1_i;
wire na770_1;
wire na770_1_i;
wire na772_2;
wire na772_2_i;
wire na774_1;
wire na774_1_i;
wire na775_1;
wire na775_1_i;
wire na775_2;
wire na775_2_i;
wire na776_1;
wire na776_1_i;
wire na776_2;
wire na776_2_i;
wire na777_1;
wire na777_1_i;
wire na777_2;
wire na777_2_i;
wire na778_1;
wire na778_1_i;
wire na778_2;
wire na778_2_i;
wire na779_1;
wire na779_1_i;
wire na779_2;
wire na779_2_i;
wire na780_1;
wire na780_1_i;
wire na780_2;
wire na780_2_i;
wire na781_1;
wire na781_1_i;
wire na781_2;
wire na781_2_i;
wire na782_1;
wire na782_1_i;
wire na782_2;
wire na782_2_i;
wire na783_1;
wire na783_1_i;
wire na783_2;
wire na783_2_i;
wire na784_1;
wire na784_1_i;
wire na784_2;
wire na784_2_i;
wire na785_1;
wire na785_1_i;
wire na785_2;
wire na785_2_i;
wire na786_1;
wire na786_1_i;
wire na786_2;
wire na786_2_i;
wire na787_1;
wire na787_1_i;
wire na787_2;
wire na787_2_i;
wire na788_1;
wire na788_1_i;
wire na788_2;
wire na788_2_i;
wire na789_1;
wire na789_1_i;
wire na789_2;
wire na789_2_i;
wire na790_1;
wire na790_1_i;
wire na790_2;
wire na790_2_i;
wire na791_1;
wire na791_1_i;
wire na791_2;
wire na791_2_i;
wire na792_1;
wire na792_1_i;
wire na792_2;
wire na792_2_i;
wire na793_1;
wire na793_1_i;
wire na793_2;
wire na793_2_i;
wire na794_1;
wire na794_1_i;
wire na794_2;
wire na794_2_i;
wire na795_1;
wire na795_1_i;
wire na795_2;
wire na795_2_i;
wire na796_1;
wire na796_1_i;
wire na796_2;
wire na796_2_i;
wire na797_1;
wire na797_1_i;
wire na797_2;
wire na797_2_i;
wire na798_1;
wire na798_1_i;
wire na798_2;
wire na798_2_i;
wire na799_1;
wire na799_1_i;
wire na799_2;
wire na799_2_i;
wire na800_1;
wire na800_1_i;
wire na800_2;
wire na800_2_i;
wire na801_1;
wire na801_1_i;
wire na801_2;
wire na801_2_i;
wire na802_1;
wire na802_1_i;
wire na802_2;
wire na802_2_i;
wire na844_2;
wire na844_2_i;
wire na862_1;
wire na862_1_i;
wire na862_2;
wire na862_2_i;
wire na866_1;
wire na866_1_i;
wire na866_2;
wire na866_2_i;
wire na868_1;
wire na868_1_i;
wire na871_1;
wire na871_1_i;
wire na871_2;
wire na871_2_i;
wire na875_2;
wire na875_2_i;
wire na876_2;
wire na876_2_i;
wire na889_1;
wire na889_1_i;
wire na889_2;
wire na889_2_i;
wire na891_1;
wire na891_1_i;
wire na891_2;
wire na891_2_i;
wire na893_1;
wire na893_1_i;
wire na893_2;
wire na893_2_i;
wire na895_1;
wire na895_1_i;
wire na895_2;
wire na895_2_i;
wire na897_1;
wire na897_1_i;
wire na897_2;
wire na897_2_i;
wire na899_1;
wire na899_1_i;
wire na899_2;
wire na899_2_i;
wire na901_1;
wire na901_1_i;
wire na901_2;
wire na901_2_i;
wire na904_2;
wire na904_2_i;
wire na906_2;
wire na906_2_i;
wire na908_1;
wire na908_1_i;
wire na925_2;
wire na925_2_i;
wire na927_2;
wire na927_2_i;
wire na929_1;
wire na929_1_i;
wire na931_1;
wire na931_1_i;
wire na933_2;
wire na933_2_i;
wire na935_2;
wire na935_2_i;
wire na937_1;
wire na937_1_i;
wire na940_2;
wire na940_2_i;
wire na941_1;
wire na941_4;
wire na942_1;
wire na942_2;
wire na942_4;
wire na944_1;
wire na944_2;
wire na944_4;
wire na946_1;
wire na946_2;
wire na948_1;
wire na949_1;
wire na949_2;
wire na949_4;
wire na951_1;
wire na951_2;
wire na951_4;
wire na953_1;
wire na953_2;
wire na953_4;
wire na955_1;
wire na955_2;
wire na955_4;
wire na957_1;
wire na957_1_i;
wire na957_2;
wire na957_4;
wire na958_1;
wire na958_1_i;
wire na958_2;
wire na958_4;
wire na960_1;
wire na960_1_i;
wire na960_2;
wire na960_4;
wire na962_1;
wire na962_1_i;
wire na962_4;
wire na963_1;
wire na963_1_i;
wire na965_1;
wire na965_1_i;
wire na965_2;
wire na965_4;
wire na967_1;
wire na967_1_i;
wire na967_2;
wire na967_4;
wire na969_1;
wire na969_1_i;
wire na969_2;
wire na969_4;
wire na971_1;
wire na971_1_i;
wire na971_2;
wire na971_4;
wire na973_1;
wire na973_1_i;
wire na973_2;
wire na973_4;
wire na974_1;
wire na974_1_i;
wire na974_2;
wire na974_4;
wire na976_1;
wire na976_1_i;
wire na976_2;
wire na976_4;
wire na978_1;
wire na978_1_i;
wire na978_4;
wire na979_1;
wire na979_1_i;
wire na981_1;
wire na981_1_i;
wire na981_2;
wire na981_4;
wire na983_1;
wire na983_1_i;
wire na983_2;
wire na983_4;
wire na985_1;
wire na985_1_i;
wire na985_2;
wire na985_4;
wire na987_1;
wire na987_1_i;
wire na987_2;
wire na987_4;
wire na989_1;
wire na990_1;
wire na990_1_i;
wire na991_1;
wire na992_1;
wire na993_1;
wire na993_1_i;
wire na994_1;
wire na995_1;
wire na996_1;
wire na996_1_i;
wire na997_1;
wire na998_1;
wire na998_1_i;
wire na999_1;
wire na1000_1;
wire na1001_1;
wire na1001_1_i;
wire na1002_1;
wire na1003_1;
wire na1004_1;
wire na1004_1_i;
wire na1005_1;
wire na1006_1;
wire na1007_1;
wire na1007_1_i;
wire na1008_1;
wire na1009_1;
wire na1009_1_i;
wire na1010_1;
wire na1011_1;
wire na1012_1;
wire na1013_1;
wire na1014_1;
wire na1015_1;
wire na1016_1;
wire na1017_1;
wire na1018_1;
wire na1019_1;
wire na1020_1;
wire na1021_1;
wire na1022_1;
wire na1023_1;
wire na1024_1;
wire na1025_1;
wire na1026_1;
wire na1027_1;
wire na1028_1;
wire na1029_2;
wire na1030_1;
wire na1032_1;
wire na1033_1;
wire na1036_1;
wire na1036_4;
wire na1037_1;
wire na1037_4;
wire na1038_3;
wire na1038_4;
wire na1038_5;
wire na1038_6;
wire na1039_3;
wire na1039_4;
wire na1039_5;
wire na1039_6;
wire na1040_1;
wire na1040_2;
wire na1041_2;
wire na1042_1;
wire na1043_2;
wire na1044_1;
wire na1045_2;
wire na1046_1;
wire na1047_2;
wire na1048_1;
wire na1049_2;
wire na1050_1;
wire na1050_4;
wire na1051_1;
wire na1052_1;
wire na1054_1;
wire na1055_2;
wire na1056_1;
wire na1060_1;
wire na1061_1;
wire na1062_1;
wire na1063_1;
wire na1064_1;
wire na1065_1;
wire na1066_1;
wire na1067_1;
wire na1068_1;
wire na1069_1;
wire na1070_1;
wire na1071_1;
wire na1072_1;
wire na1073_1;
wire na1075_1;
wire na1076_2;
wire na1079_1;
wire na1080_1;
wire na1081_1;
wire na1082_1;
wire na1083_1;
wire na1084_1;
wire na1085_1;
wire na1087_1;
wire na1088_1;
wire na1090_2;
wire na1091_1;
wire na1092_1;
wire na1092_2;
wire na1095_1;
wire na1095_2;
wire na1097_1;
wire na1098_1;
wire na1098_2;
wire na1100_1;
wire na1102_2;
wire na1112_1;
wire na1112_2;
wire na1113_2;
wire na1114_1;
wire na1114_2;
wire na1116_1;
wire na1118_2;
wire na1128_1;
wire na1128_2;
wire na1129_1;
wire na1130_2;
wire na1131_1;
wire na1131_2;
wire na1131_3;
wire na1131_3_i;
wire na1131_6;
wire na1132_1;
wire na1132_1_i;
wire na1132_2;
wire na1132_2_i;
wire na1132_3;
wire na1132_6;
wire na1133_1;
wire na1133_1_i;
wire na1133_2;
wire na1133_2_i;
wire na1133_3;
wire na1133_6;
wire na1134_1;
wire na1134_1_i;
wire na1134_2;
wire na1134_2_i;
wire na1134_3;
wire na1134_6;
wire na1135_1;
wire na1135_1_i;
wire na1135_2;
wire na1135_2_i;
wire na1135_3;
wire na1135_6;
wire na1136_1;
wire na1136_1_i;
wire na1136_2;
wire na1136_2_i;
wire na1136_3;
wire na1136_6;
wire na1137_1;
wire na1137_1_i;
wire na1137_2;
wire na1137_2_i;
wire na1137_3;
wire na1137_6;
wire na1138_1;
wire na1138_1_i;
wire na1138_2;
wire na1138_2_i;
wire na1138_3;
wire na1138_6;
wire na1139_1;
wire na1139_1_i;
wire na1139_2;
wire na1139_2_i;
wire na1139_3;
wire na1139_6;
wire na1140_1;
wire na1140_1_i;
wire na1140_2;
wire na1140_2_i;
wire na1140_3;
wire na1140_6;
wire na1141_1;
wire na1141_1_i;
wire na1141_2;
wire na1141_2_i;
wire na1141_3;
wire na1141_6;
wire na1142_1;
wire na1142_1_i;
wire na1142_2;
wire na1142_2_i;
wire na1142_3;
wire na1142_6;
wire na1143_1;
wire na1143_1_i;
wire na1143_2;
wire na1143_2_i;
wire na1143_3;
wire na1143_6;
wire na1144_1;
wire na1144_1_i;
wire na1144_2;
wire na1144_2_i;
wire na1144_3;
wire na1144_6;
wire na1145_1;
wire na1145_1_i;
wire na1145_2;
wire na1145_2_i;
wire na1145_3;
wire na1145_6;
wire na1146_1;
wire na1146_1_i;
wire na1146_2;
wire na1146_2_i;
wire na1146_3;
wire na1146_6;
wire na1147_1;
wire na1147_1_i;
wire na1147_2;
wire na1147_2_i;
wire na1147_3;
wire na1147_6;
wire na1148_1;
wire na1148_2;
wire na1148_4;
wire na1148_7;
wire na1149_1;
wire na1149_3_i;
wire na1149_4;
wire na1149_5;
wire na1149_7;
wire na1150_3;
wire na1150_4;
wire na1150_5;
wire na1150_7;
wire na1151_1;
wire na1151_2;
wire na1151_3;
wire na1151_3_i;
wire na1151_4;
wire na1151_5;
wire na1151_7;
wire na1151_8;
wire na1152_4;
wire na1152_5;
wire na1152_7;
wire na1152_8;
wire na1153_3;
wire na1153_4;
wire na1153_5;
wire na1153_6;
wire na1153_7;
wire na1153_8;
wire na1154_3;
wire na1154_4;
wire na1154_5;
wire na1154_6;
wire na1154_7;
wire na1154_8;
wire na1155_3;
wire na1155_4;
wire na1155_5;
wire na1155_6;
wire na1155_7;
wire na1155_8;
wire na1156_3;
wire na1156_4;
wire na1156_5;
wire na1156_6;
wire na1156_7;
wire na1156_8;
wire na1157_3;
wire na1157_4;
wire na1157_5;
wire na1157_6;
wire na1157_7;
wire na1157_8;
wire na1158_3;
wire na1158_4;
wire na1158_5;
wire na1158_6;
wire na1158_7;
wire na1158_8;
wire na1159_3;
wire na1159_4;
wire na1159_5;
wire na1159_6;
wire na1159_7;
wire na1159_8;
wire na1160_3;
wire na1160_4;
wire na1160_5;
wire na1160_6;
wire na1160_7;
wire na1160_8;
wire na1161_3;
wire na1161_4;
wire na1161_5;
wire na1161_6;
wire na1161_7;
wire na1161_8;
wire na1162_3;
wire na1162_4;
wire na1162_5;
wire na1162_6;
wire na1162_7;
wire na1162_8;
wire na1163_3;
wire na1163_4;
wire na1163_5;
wire na1163_6;
wire na1163_7;
wire na1163_8;
wire na1164_3;
wire na1164_4;
wire na1164_5;
wire na1164_6;
wire na1164_7;
wire na1164_8;
wire na1165_3;
wire na1165_4;
wire na1165_5;
wire na1165_6;
wire na1165_7;
wire na1165_8;
wire na1166_3;
wire na1166_4;
wire na1166_5;
wire na1166_6;
wire na1166_7;
wire na1166_8;
wire na1167_3;
wire na1167_4;
wire na1167_5;
wire na1167_6;
wire na1167_7;
wire na1167_8;
wire na1168_3;
wire na1168_4;
wire na1168_5;
wire na1168_6;
wire na1168_7;
wire na1168_8;
wire na1169_2;
wire na1169_3;
wire na1169_3_i;
wire na1169_6;
wire na1170_1;
wire na1170_2;
wire na1170_4;
wire na1170_7;
wire na1171_1;
wire na1171_3_i;
wire na1171_4;
wire na1171_5;
wire na1171_7;
wire na1172_3;
wire na1172_4;
wire na1172_5;
wire na1172_7;
wire na1173_1;
wire na1173_2;
wire na1173_3;
wire na1173_3_i;
wire na1173_4;
wire na1173_5;
wire na1173_7;
wire na1173_8;
wire na1174_4;
wire na1174_5;
wire na1174_7;
wire na1174_8;
wire na1175_3;
wire na1175_4;
wire na1175_5;
wire na1175_6;
wire na1175_7;
wire na1175_8;
wire na1176_3;
wire na1176_4;
wire na1176_5;
wire na1176_6;
wire na1176_7;
wire na1176_8;
wire na1177_3;
wire na1177_4;
wire na1177_5;
wire na1177_6;
wire na1177_7;
wire na1177_8;
wire na1178_3;
wire na1178_4;
wire na1178_5;
wire na1178_6;
wire na1178_7;
wire na1178_8;
wire na1179_3;
wire na1179_4;
wire na1179_5;
wire na1179_6;
wire na1179_7;
wire na1179_8;
wire na1180_3;
wire na1180_4;
wire na1180_5;
wire na1180_6;
wire na1180_7;
wire na1180_8;
wire na1181_3;
wire na1181_4;
wire na1181_5;
wire na1181_6;
wire na1181_7;
wire na1181_8;
wire na1182_3;
wire na1182_4;
wire na1182_5;
wire na1182_6;
wire na1182_7;
wire na1182_8;
wire na1183_3;
wire na1183_4;
wire na1183_5;
wire na1183_6;
wire na1183_7;
wire na1183_8;
wire na1184_3;
wire na1184_4;
wire na1184_5;
wire na1184_6;
wire na1184_7;
wire na1184_8;
wire na1185_3;
wire na1185_4;
wire na1185_5;
wire na1185_6;
wire na1185_7;
wire na1185_8;
wire na1186_3;
wire na1186_4;
wire na1186_5;
wire na1186_6;
wire na1186_7;
wire na1186_8;
wire na1187_3;
wire na1187_4;
wire na1187_5;
wire na1187_6;
wire na1187_7;
wire na1187_8;
wire na1188_3;
wire na1188_4;
wire na1188_5;
wire na1188_6;
wire na1188_7;
wire na1188_8;
wire na1189_3;
wire na1189_4;
wire na1189_5;
wire na1189_6;
wire na1189_7;
wire na1189_8;
wire na1190_3;
wire na1190_4;
wire na1190_5;
wire na1190_6;
wire na1190_7;
wire na1190_8;
wire na1191_2;
wire na1191_3;
wire na1191_3_i;
wire na1191_6;
wire na1192_1;
wire na1192_2;
wire na1192_4;
wire na1192_7;
wire na1193_1;
wire na1193_3_i;
wire na1193_4;
wire na1193_5;
wire na1193_7;
wire na1194_3;
wire na1194_4;
wire na1194_5;
wire na1194_7;
wire na1195_1;
wire na1195_2;
wire na1195_3;
wire na1195_3_i;
wire na1195_4;
wire na1195_5;
wire na1195_7;
wire na1195_8;
wire na1196_4;
wire na1196_5;
wire na1196_7;
wire na1196_8;
wire na1197_3;
wire na1197_4;
wire na1197_5;
wire na1197_6;
wire na1197_7;
wire na1197_8;
wire na1198_3;
wire na1198_4;
wire na1198_5;
wire na1198_6;
wire na1198_7;
wire na1198_8;
wire na1199_3;
wire na1199_4;
wire na1199_5;
wire na1199_6;
wire na1199_7;
wire na1199_8;
wire na1200_3;
wire na1200_4;
wire na1200_5;
wire na1200_6;
wire na1200_7;
wire na1200_8;
wire na1201_3;
wire na1201_4;
wire na1201_5;
wire na1201_6;
wire na1201_7;
wire na1201_8;
wire na1202_3;
wire na1202_4;
wire na1202_5;
wire na1202_6;
wire na1202_7;
wire na1202_8;
wire na1203_3;
wire na1203_4;
wire na1203_5;
wire na1203_6;
wire na1203_7;
wire na1203_8;
wire na1204_3;
wire na1204_4;
wire na1204_5;
wire na1204_6;
wire na1204_7;
wire na1204_8;
wire na1205_3;
wire na1205_4;
wire na1205_5;
wire na1205_6;
wire na1205_7;
wire na1205_8;
wire na1206_3;
wire na1206_4;
wire na1206_5;
wire na1206_6;
wire na1206_7;
wire na1206_8;
wire na1207_3;
wire na1207_4;
wire na1207_5;
wire na1207_6;
wire na1207_7;
wire na1207_8;
wire na1208_3;
wire na1208_4;
wire na1208_5;
wire na1208_6;
wire na1208_7;
wire na1208_8;
wire na1209_3;
wire na1209_4;
wire na1209_5;
wire na1209_6;
wire na1209_7;
wire na1209_8;
wire na1210_3;
wire na1210_4;
wire na1210_5;
wire na1210_6;
wire na1210_7;
wire na1210_8;
wire na1211_3;
wire na1211_4;
wire na1211_5;
wire na1211_6;
wire na1211_7;
wire na1211_8;
wire na1212_3;
wire na1212_4;
wire na1212_5;
wire na1212_6;
wire na1212_7;
wire na1212_8;
wire na1213_2;
wire na1213_3;
wire na1213_3_i;
wire na1213_6;
wire na1214_1;
wire na1214_2;
wire na1214_4;
wire na1214_7;
wire na1215_1;
wire na1215_3_i;
wire na1215_4;
wire na1215_5;
wire na1215_7;
wire na1216_3;
wire na1216_4;
wire na1216_5;
wire na1216_7;
wire na1217_1;
wire na1217_2;
wire na1217_3;
wire na1217_3_i;
wire na1217_4;
wire na1217_5;
wire na1217_7;
wire na1217_8;
wire na1218_4;
wire na1218_5;
wire na1218_7;
wire na1218_8;
wire na1219_3;
wire na1219_4;
wire na1219_5;
wire na1219_6;
wire na1219_7;
wire na1219_8;
wire na1220_3;
wire na1220_4;
wire na1220_5;
wire na1220_6;
wire na1220_7;
wire na1220_8;
wire na1221_3;
wire na1221_4;
wire na1221_5;
wire na1221_6;
wire na1221_7;
wire na1221_8;
wire na1222_3;
wire na1222_4;
wire na1222_5;
wire na1222_6;
wire na1222_7;
wire na1222_8;
wire na1223_3;
wire na1223_4;
wire na1223_5;
wire na1223_6;
wire na1223_7;
wire na1223_8;
wire na1224_3;
wire na1224_4;
wire na1224_5;
wire na1224_6;
wire na1224_7;
wire na1224_8;
wire na1225_3;
wire na1225_4;
wire na1225_5;
wire na1225_6;
wire na1225_7;
wire na1225_8;
wire na1226_3;
wire na1226_4;
wire na1226_5;
wire na1226_6;
wire na1226_7;
wire na1226_8;
wire na1227_3;
wire na1227_4;
wire na1227_5;
wire na1227_6;
wire na1227_7;
wire na1227_8;
wire na1228_3;
wire na1228_4;
wire na1228_5;
wire na1228_6;
wire na1228_7;
wire na1228_8;
wire na1229_3;
wire na1229_4;
wire na1229_5;
wire na1229_6;
wire na1229_7;
wire na1229_8;
wire na1230_3;
wire na1230_4;
wire na1230_5;
wire na1230_6;
wire na1230_7;
wire na1230_8;
wire na1231_3;
wire na1231_4;
wire na1231_5;
wire na1231_6;
wire na1231_7;
wire na1231_8;
wire na1232_3;
wire na1232_4;
wire na1232_5;
wire na1232_6;
wire na1232_7;
wire na1232_8;
wire na1233_3;
wire na1233_4;
wire na1233_5;
wire na1233_6;
wire na1233_7;
wire na1233_8;
wire na1234_3;
wire na1234_4;
wire na1234_5;
wire na1234_6;
wire na1234_7;
wire na1234_8;
wire na1235_2;
wire na1235_3;
wire na1235_3_i;
wire na1235_6;
wire na1236_1;
wire na1236_2;
wire na1236_4;
wire na1236_7;
wire na1237_1;
wire na1237_3_i;
wire na1237_4;
wire na1237_5;
wire na1237_7;
wire na1238_3;
wire na1238_4;
wire na1238_5;
wire na1238_7;
wire na1239_1;
wire na1239_2;
wire na1239_3;
wire na1239_3_i;
wire na1239_4;
wire na1239_5;
wire na1239_7;
wire na1239_8;
wire na1240_4;
wire na1240_5;
wire na1240_7;
wire na1240_8;
wire na1241_3;
wire na1241_4;
wire na1241_5;
wire na1241_6;
wire na1241_7;
wire na1241_8;
wire na1242_3;
wire na1242_4;
wire na1242_5;
wire na1242_6;
wire na1242_7;
wire na1242_8;
wire na1243_3;
wire na1243_4;
wire na1243_5;
wire na1243_6;
wire na1243_7;
wire na1243_8;
wire na1244_3;
wire na1244_4;
wire na1244_5;
wire na1244_6;
wire na1244_7;
wire na1244_8;
wire na1245_3;
wire na1245_4;
wire na1245_5;
wire na1245_6;
wire na1245_7;
wire na1245_8;
wire na1246_3;
wire na1246_4;
wire na1246_5;
wire na1246_6;
wire na1246_7;
wire na1246_8;
wire na1247_3;
wire na1247_4;
wire na1247_5;
wire na1247_6;
wire na1247_7;
wire na1247_8;
wire na1248_3;
wire na1248_4;
wire na1248_5;
wire na1248_6;
wire na1248_7;
wire na1248_8;
wire na1249_3;
wire na1249_4;
wire na1249_5;
wire na1249_6;
wire na1249_7;
wire na1249_8;
wire na1250_3;
wire na1250_4;
wire na1250_5;
wire na1250_6;
wire na1250_7;
wire na1250_8;
wire na1251_3;
wire na1251_4;
wire na1251_5;
wire na1251_6;
wire na1251_7;
wire na1251_8;
wire na1252_3;
wire na1252_4;
wire na1252_5;
wire na1252_6;
wire na1252_7;
wire na1252_8;
wire na1253_3;
wire na1253_4;
wire na1253_5;
wire na1253_6;
wire na1253_7;
wire na1253_8;
wire na1254_3;
wire na1254_4;
wire na1254_5;
wire na1254_6;
wire na1254_7;
wire na1254_8;
wire na1255_3;
wire na1255_4;
wire na1255_5;
wire na1255_6;
wire na1255_7;
wire na1255_8;
wire na1256_3;
wire na1256_4;
wire na1256_5;
wire na1256_6;
wire na1256_7;
wire na1256_8;
wire na1257_2;
wire na1257_3;
wire na1257_3_i;
wire na1257_6;
wire na1258_1;
wire na1258_2;
wire na1258_4;
wire na1258_7;
wire na1259_1;
wire na1259_3_i;
wire na1259_4;
wire na1259_5;
wire na1259_7;
wire na1260_3;
wire na1260_4;
wire na1260_5;
wire na1260_7;
wire na1261_1;
wire na1261_2;
wire na1261_3;
wire na1261_3_i;
wire na1261_4;
wire na1261_5;
wire na1261_7;
wire na1261_8;
wire na1262_4;
wire na1262_5;
wire na1262_7;
wire na1262_8;
wire na1263_3;
wire na1263_4;
wire na1263_5;
wire na1263_6;
wire na1263_7;
wire na1263_8;
wire na1264_3;
wire na1264_4;
wire na1264_5;
wire na1264_6;
wire na1264_7;
wire na1264_8;
wire na1265_3;
wire na1265_4;
wire na1265_5;
wire na1265_6;
wire na1265_7;
wire na1265_8;
wire na1266_3;
wire na1266_4;
wire na1266_5;
wire na1266_6;
wire na1266_7;
wire na1266_8;
wire na1267_3;
wire na1267_4;
wire na1267_5;
wire na1267_6;
wire na1267_7;
wire na1267_8;
wire na1268_3;
wire na1268_4;
wire na1268_5;
wire na1268_6;
wire na1268_7;
wire na1268_8;
wire na1269_3;
wire na1269_4;
wire na1269_5;
wire na1269_6;
wire na1269_7;
wire na1269_8;
wire na1270_3;
wire na1270_4;
wire na1270_5;
wire na1270_6;
wire na1270_7;
wire na1270_8;
wire na1271_3;
wire na1271_4;
wire na1271_5;
wire na1271_6;
wire na1271_7;
wire na1271_8;
wire na1272_3;
wire na1272_4;
wire na1272_5;
wire na1272_6;
wire na1272_7;
wire na1272_8;
wire na1273_3;
wire na1273_4;
wire na1273_5;
wire na1273_6;
wire na1273_7;
wire na1273_8;
wire na1274_3;
wire na1274_4;
wire na1274_5;
wire na1274_6;
wire na1274_7;
wire na1274_8;
wire na1275_3;
wire na1275_4;
wire na1275_5;
wire na1275_6;
wire na1275_7;
wire na1275_8;
wire na1276_3;
wire na1276_4;
wire na1276_5;
wire na1276_6;
wire na1276_7;
wire na1276_8;
wire na1277_3;
wire na1277_4;
wire na1277_5;
wire na1277_6;
wire na1277_7;
wire na1277_8;
wire na1278_3;
wire na1278_4;
wire na1278_5;
wire na1278_6;
wire na1278_7;
wire na1278_8;
wire na1279_2;
wire na1279_3;
wire na1279_3_i;
wire na1279_6;
wire na1280_1;
wire na1280_2;
wire na1280_4;
wire na1280_7;
wire na1281_1;
wire na1281_3_i;
wire na1281_4;
wire na1281_5;
wire na1281_7;
wire na1282_3;
wire na1282_4;
wire na1282_5;
wire na1282_7;
wire na1283_1;
wire na1283_2;
wire na1283_3;
wire na1283_3_i;
wire na1283_4;
wire na1283_5;
wire na1283_7;
wire na1283_8;
wire na1284_4;
wire na1284_5;
wire na1284_7;
wire na1284_8;
wire na1285_3;
wire na1285_4;
wire na1285_5;
wire na1285_6;
wire na1285_7;
wire na1285_8;
wire na1286_3;
wire na1286_4;
wire na1286_5;
wire na1286_6;
wire na1286_7;
wire na1286_8;
wire na1287_3;
wire na1287_4;
wire na1287_5;
wire na1287_6;
wire na1287_7;
wire na1287_8;
wire na1288_3;
wire na1288_4;
wire na1288_5;
wire na1288_6;
wire na1288_7;
wire na1288_8;
wire na1289_3;
wire na1289_4;
wire na1289_5;
wire na1289_6;
wire na1289_7;
wire na1289_8;
wire na1290_3;
wire na1290_4;
wire na1290_5;
wire na1290_6;
wire na1290_7;
wire na1290_8;
wire na1291_3;
wire na1291_4;
wire na1291_5;
wire na1291_6;
wire na1291_7;
wire na1291_8;
wire na1292_3;
wire na1292_4;
wire na1292_5;
wire na1292_6;
wire na1292_7;
wire na1292_8;
wire na1293_3;
wire na1293_4;
wire na1293_5;
wire na1293_6;
wire na1293_7;
wire na1293_8;
wire na1294_3;
wire na1294_4;
wire na1294_5;
wire na1294_6;
wire na1294_7;
wire na1294_8;
wire na1295_3;
wire na1295_4;
wire na1295_5;
wire na1295_6;
wire na1295_7;
wire na1295_8;
wire na1296_3;
wire na1296_4;
wire na1296_5;
wire na1296_6;
wire na1296_7;
wire na1296_8;
wire na1297_3;
wire na1297_4;
wire na1297_5;
wire na1297_6;
wire na1297_7;
wire na1297_8;
wire na1298_3;
wire na1298_4;
wire na1298_5;
wire na1298_6;
wire na1298_7;
wire na1298_8;
wire na1299_3;
wire na1299_4;
wire na1299_5;
wire na1299_6;
wire na1299_7;
wire na1299_8;
wire na1300_3;
wire na1300_4;
wire na1300_5;
wire na1300_6;
wire na1300_7;
wire na1300_8;
wire na1301_2;
wire na1301_3;
wire na1301_3_i;
wire na1301_6;
wire na1302_1;
wire na1302_2;
wire na1302_4;
wire na1302_7;
wire na1303_1;
wire na1303_3_i;
wire na1303_4;
wire na1303_5;
wire na1303_7;
wire na1304_3;
wire na1304_4;
wire na1304_5;
wire na1304_7;
wire na1305_1;
wire na1305_2;
wire na1305_3;
wire na1305_3_i;
wire na1305_4;
wire na1305_5;
wire na1305_7;
wire na1305_8;
wire na1306_4;
wire na1306_5;
wire na1306_7;
wire na1306_8;
wire na1307_3;
wire na1307_4;
wire na1307_5;
wire na1307_6;
wire na1307_7;
wire na1307_8;
wire na1308_3;
wire na1308_4;
wire na1308_5;
wire na1308_6;
wire na1308_7;
wire na1308_8;
wire na1309_3;
wire na1309_4;
wire na1309_5;
wire na1309_6;
wire na1309_7;
wire na1309_8;
wire na1310_3;
wire na1310_4;
wire na1310_5;
wire na1310_6;
wire na1310_7;
wire na1310_8;
wire na1311_3;
wire na1311_4;
wire na1311_5;
wire na1311_6;
wire na1311_7;
wire na1311_8;
wire na1312_3;
wire na1312_4;
wire na1312_5;
wire na1312_6;
wire na1312_7;
wire na1312_8;
wire na1313_3;
wire na1313_4;
wire na1313_5;
wire na1313_6;
wire na1313_7;
wire na1313_8;
wire na1314_3;
wire na1314_4;
wire na1314_5;
wire na1314_6;
wire na1314_7;
wire na1314_8;
wire na1315_3;
wire na1315_4;
wire na1315_5;
wire na1315_6;
wire na1315_7;
wire na1315_8;
wire na1316_3;
wire na1316_4;
wire na1316_5;
wire na1316_6;
wire na1316_7;
wire na1316_8;
wire na1317_3;
wire na1317_4;
wire na1317_5;
wire na1317_6;
wire na1317_7;
wire na1317_8;
wire na1318_3;
wire na1318_4;
wire na1318_5;
wire na1318_6;
wire na1318_7;
wire na1318_8;
wire na1319_3;
wire na1319_4;
wire na1319_5;
wire na1319_6;
wire na1319_7;
wire na1319_8;
wire na1320_3;
wire na1320_4;
wire na1320_5;
wire na1320_6;
wire na1320_7;
wire na1320_8;
wire na1321_3;
wire na1321_4;
wire na1321_5;
wire na1321_6;
wire na1321_7;
wire na1321_8;
wire na1322_3;
wire na1322_4;
wire na1322_5;
wire na1322_6;
wire na1322_7;
wire na1322_8;
wire na1323_2;
wire na1323_3;
wire na1323_3_i;
wire na1323_6;
wire na1324_1;
wire na1324_2;
wire na1324_4;
wire na1324_7;
wire na1325_1;
wire na1325_3_i;
wire na1325_4;
wire na1325_5;
wire na1325_7;
wire na1326_3;
wire na1326_4;
wire na1326_5;
wire na1326_7;
wire na1327_1;
wire na1327_2;
wire na1327_3;
wire na1327_3_i;
wire na1327_4;
wire na1327_5;
wire na1327_7;
wire na1327_8;
wire na1328_4;
wire na1328_5;
wire na1328_7;
wire na1328_8;
wire na1329_3;
wire na1329_4;
wire na1329_5;
wire na1329_6;
wire na1329_7;
wire na1329_8;
wire na1330_3;
wire na1330_4;
wire na1330_5;
wire na1330_6;
wire na1330_7;
wire na1330_8;
wire na1331_3;
wire na1331_4;
wire na1331_5;
wire na1331_6;
wire na1331_7;
wire na1331_8;
wire na1332_3;
wire na1332_4;
wire na1332_5;
wire na1332_6;
wire na1332_7;
wire na1332_8;
wire na1333_3;
wire na1333_4;
wire na1333_5;
wire na1333_6;
wire na1333_7;
wire na1333_8;
wire na1334_3;
wire na1334_4;
wire na1334_5;
wire na1334_6;
wire na1334_7;
wire na1334_8;
wire na1335_3;
wire na1335_4;
wire na1335_5;
wire na1335_6;
wire na1335_7;
wire na1335_8;
wire na1336_3;
wire na1336_4;
wire na1336_5;
wire na1336_6;
wire na1336_7;
wire na1336_8;
wire na1337_3;
wire na1337_4;
wire na1337_5;
wire na1337_6;
wire na1337_7;
wire na1337_8;
wire na1338_3;
wire na1338_4;
wire na1338_5;
wire na1338_6;
wire na1338_7;
wire na1338_8;
wire na1339_3;
wire na1339_4;
wire na1339_5;
wire na1339_6;
wire na1339_7;
wire na1339_8;
wire na1340_3;
wire na1340_4;
wire na1340_5;
wire na1340_6;
wire na1340_7;
wire na1340_8;
wire na1341_3;
wire na1341_4;
wire na1341_5;
wire na1341_6;
wire na1341_7;
wire na1341_8;
wire na1342_3;
wire na1342_4;
wire na1342_5;
wire na1342_6;
wire na1342_7;
wire na1342_8;
wire na1343_3;
wire na1343_4;
wire na1343_5;
wire na1343_6;
wire na1343_7;
wire na1343_8;
wire na1344_3;
wire na1344_4;
wire na1344_5;
wire na1344_6;
wire na1344_7;
wire na1344_8;
wire na1345_2;
wire na1345_3;
wire na1345_3_i;
wire na1345_6;
wire na1346_1;
wire na1346_2;
wire na1346_4;
wire na1346_7;
wire na1347_1;
wire na1347_3_i;
wire na1347_4;
wire na1347_5;
wire na1347_7;
wire na1348_3;
wire na1348_4;
wire na1348_5;
wire na1348_7;
wire na1349_1;
wire na1349_2;
wire na1349_3;
wire na1349_3_i;
wire na1349_4;
wire na1349_5;
wire na1349_7;
wire na1349_8;
wire na1350_4;
wire na1350_5;
wire na1350_7;
wire na1350_8;
wire na1351_3;
wire na1351_4;
wire na1351_5;
wire na1351_6;
wire na1351_7;
wire na1351_8;
wire na1352_3;
wire na1352_4;
wire na1352_5;
wire na1352_6;
wire na1352_7;
wire na1352_8;
wire na1353_3;
wire na1353_4;
wire na1353_5;
wire na1353_6;
wire na1353_7;
wire na1353_8;
wire na1354_3;
wire na1354_4;
wire na1354_5;
wire na1354_6;
wire na1354_7;
wire na1354_8;
wire na1355_3;
wire na1355_4;
wire na1355_5;
wire na1355_6;
wire na1355_7;
wire na1355_8;
wire na1356_3;
wire na1356_4;
wire na1356_5;
wire na1356_6;
wire na1356_7;
wire na1356_8;
wire na1357_3;
wire na1357_4;
wire na1357_5;
wire na1357_6;
wire na1357_7;
wire na1357_8;
wire na1358_3;
wire na1358_4;
wire na1358_5;
wire na1358_6;
wire na1358_7;
wire na1358_8;
wire na1359_3;
wire na1359_4;
wire na1359_5;
wire na1359_6;
wire na1359_7;
wire na1359_8;
wire na1360_3;
wire na1360_4;
wire na1360_5;
wire na1360_6;
wire na1360_7;
wire na1360_8;
wire na1361_3;
wire na1361_4;
wire na1361_5;
wire na1361_6;
wire na1361_7;
wire na1361_8;
wire na1362_3;
wire na1362_4;
wire na1362_5;
wire na1362_6;
wire na1362_7;
wire na1362_8;
wire na1363_3;
wire na1363_4;
wire na1363_5;
wire na1363_6;
wire na1363_7;
wire na1363_8;
wire na1364_3;
wire na1364_4;
wire na1364_5;
wire na1364_6;
wire na1364_7;
wire na1364_8;
wire na1365_3;
wire na1365_4;
wire na1365_5;
wire na1365_6;
wire na1365_7;
wire na1365_8;
wire na1366_3;
wire na1366_4;
wire na1366_5;
wire na1366_6;
wire na1366_7;
wire na1366_8;
wire na1367_2;
wire na1367_3;
wire na1367_3_i;
wire na1367_6;
wire na1368_1;
wire na1368_2;
wire na1368_4;
wire na1368_7;
wire na1369_1;
wire na1369_3_i;
wire na1369_4;
wire na1369_5;
wire na1369_7;
wire na1370_3;
wire na1370_4;
wire na1370_5;
wire na1370_7;
wire na1371_1;
wire na1371_2;
wire na1371_3;
wire na1371_3_i;
wire na1371_4;
wire na1371_5;
wire na1371_7;
wire na1371_8;
wire na1372_4;
wire na1372_5;
wire na1372_7;
wire na1372_8;
wire na1373_3;
wire na1373_4;
wire na1373_5;
wire na1373_6;
wire na1373_7;
wire na1373_8;
wire na1374_3;
wire na1374_4;
wire na1374_5;
wire na1374_6;
wire na1374_7;
wire na1374_8;
wire na1375_3;
wire na1375_4;
wire na1375_5;
wire na1375_6;
wire na1375_7;
wire na1375_8;
wire na1376_3;
wire na1376_4;
wire na1376_5;
wire na1376_6;
wire na1376_7;
wire na1376_8;
wire na1377_3;
wire na1377_4;
wire na1377_5;
wire na1377_6;
wire na1377_7;
wire na1377_8;
wire na1378_3;
wire na1378_4;
wire na1378_5;
wire na1378_6;
wire na1378_7;
wire na1378_8;
wire na1379_3;
wire na1379_4;
wire na1379_5;
wire na1379_6;
wire na1379_7;
wire na1379_8;
wire na1380_3;
wire na1380_4;
wire na1380_5;
wire na1380_6;
wire na1380_7;
wire na1380_8;
wire na1381_3;
wire na1381_4;
wire na1381_5;
wire na1381_6;
wire na1381_7;
wire na1381_8;
wire na1382_3;
wire na1382_4;
wire na1382_5;
wire na1382_6;
wire na1382_7;
wire na1382_8;
wire na1383_3;
wire na1383_4;
wire na1383_5;
wire na1383_6;
wire na1383_7;
wire na1383_8;
wire na1384_3;
wire na1384_4;
wire na1384_5;
wire na1384_6;
wire na1384_7;
wire na1384_8;
wire na1385_3;
wire na1385_4;
wire na1385_5;
wire na1385_6;
wire na1385_7;
wire na1385_8;
wire na1386_3;
wire na1386_4;
wire na1386_5;
wire na1386_6;
wire na1386_7;
wire na1386_8;
wire na1387_3;
wire na1387_4;
wire na1387_5;
wire na1387_6;
wire na1387_7;
wire na1387_8;
wire na1388_3;
wire na1388_4;
wire na1388_5;
wire na1388_6;
wire na1388_7;
wire na1388_8;
wire na1389_2;
wire na1389_3;
wire na1389_3_i;
wire na1389_6;
wire na1390_1;
wire na1390_2;
wire na1390_4;
wire na1390_7;
wire na1391_1;
wire na1391_3_i;
wire na1391_4;
wire na1391_5;
wire na1391_7;
wire na1392_3;
wire na1392_4;
wire na1392_5;
wire na1392_7;
wire na1393_1;
wire na1393_2;
wire na1393_3;
wire na1393_3_i;
wire na1393_4;
wire na1393_5;
wire na1393_7;
wire na1393_8;
wire na1394_4;
wire na1394_5;
wire na1394_7;
wire na1394_8;
wire na1395_3;
wire na1395_4;
wire na1395_5;
wire na1395_6;
wire na1395_7;
wire na1395_8;
wire na1396_3;
wire na1396_4;
wire na1396_5;
wire na1396_6;
wire na1396_7;
wire na1396_8;
wire na1397_3;
wire na1397_4;
wire na1397_5;
wire na1397_6;
wire na1397_7;
wire na1397_8;
wire na1398_3;
wire na1398_4;
wire na1398_5;
wire na1398_6;
wire na1398_7;
wire na1398_8;
wire na1399_3;
wire na1399_4;
wire na1399_5;
wire na1399_6;
wire na1399_7;
wire na1399_8;
wire na1400_3;
wire na1400_4;
wire na1400_5;
wire na1400_6;
wire na1400_7;
wire na1400_8;
wire na1401_3;
wire na1401_4;
wire na1401_5;
wire na1401_6;
wire na1401_7;
wire na1401_8;
wire na1402_3;
wire na1402_4;
wire na1402_5;
wire na1402_6;
wire na1402_7;
wire na1402_8;
wire na1403_3;
wire na1403_4;
wire na1403_5;
wire na1403_6;
wire na1403_7;
wire na1403_8;
wire na1404_3;
wire na1404_4;
wire na1404_5;
wire na1404_6;
wire na1404_7;
wire na1404_8;
wire na1405_3;
wire na1405_4;
wire na1405_5;
wire na1405_6;
wire na1405_7;
wire na1405_8;
wire na1406_3;
wire na1406_4;
wire na1406_5;
wire na1406_6;
wire na1406_7;
wire na1406_8;
wire na1407_3;
wire na1407_4;
wire na1407_5;
wire na1407_6;
wire na1407_7;
wire na1407_8;
wire na1408_3;
wire na1408_4;
wire na1408_5;
wire na1408_6;
wire na1408_7;
wire na1408_8;
wire na1409_3;
wire na1409_4;
wire na1409_5;
wire na1409_6;
wire na1409_7;
wire na1409_8;
wire na1410_3;
wire na1410_4;
wire na1410_5;
wire na1410_6;
wire na1410_7;
wire na1410_8;
wire na1411_2;
wire na1411_3;
wire na1411_3_i;
wire na1411_6;
wire na1412_1;
wire na1412_2;
wire na1412_4;
wire na1412_7;
wire na1413_1;
wire na1413_3_i;
wire na1413_4;
wire na1413_5;
wire na1413_7;
wire na1414_3;
wire na1414_4;
wire na1414_5;
wire na1414_7;
wire na1415_1;
wire na1415_2;
wire na1415_3;
wire na1415_3_i;
wire na1415_4;
wire na1415_5;
wire na1415_7;
wire na1415_8;
wire na1416_4;
wire na1416_5;
wire na1416_7;
wire na1416_8;
wire na1417_3;
wire na1417_4;
wire na1417_5;
wire na1417_6;
wire na1417_7;
wire na1417_8;
wire na1418_3;
wire na1418_4;
wire na1418_5;
wire na1418_6;
wire na1418_7;
wire na1418_8;
wire na1419_3;
wire na1419_4;
wire na1419_5;
wire na1419_6;
wire na1419_7;
wire na1419_8;
wire na1420_3;
wire na1420_4;
wire na1420_5;
wire na1420_6;
wire na1420_7;
wire na1420_8;
wire na1421_3;
wire na1421_4;
wire na1421_5;
wire na1421_6;
wire na1421_7;
wire na1421_8;
wire na1422_3;
wire na1422_4;
wire na1422_5;
wire na1422_6;
wire na1422_7;
wire na1422_8;
wire na1423_3;
wire na1423_4;
wire na1423_5;
wire na1423_6;
wire na1423_7;
wire na1423_8;
wire na1424_3;
wire na1424_4;
wire na1424_5;
wire na1424_6;
wire na1424_7;
wire na1424_8;
wire na1425_3;
wire na1425_4;
wire na1425_5;
wire na1425_6;
wire na1425_7;
wire na1425_8;
wire na1426_3;
wire na1426_4;
wire na1426_5;
wire na1426_6;
wire na1426_7;
wire na1426_8;
wire na1427_3;
wire na1427_4;
wire na1427_5;
wire na1427_6;
wire na1427_7;
wire na1427_8;
wire na1428_3;
wire na1428_4;
wire na1428_5;
wire na1428_6;
wire na1428_7;
wire na1428_8;
wire na1429_3;
wire na1429_4;
wire na1429_5;
wire na1429_6;
wire na1429_7;
wire na1429_8;
wire na1430_3;
wire na1430_4;
wire na1430_5;
wire na1430_6;
wire na1430_7;
wire na1430_8;
wire na1431_3;
wire na1431_4;
wire na1431_5;
wire na1431_6;
wire na1431_7;
wire na1431_8;
wire na1432_3;
wire na1432_4;
wire na1432_5;
wire na1432_6;
wire na1432_7;
wire na1432_8;
wire na1433_2;
wire na1433_3;
wire na1433_3_i;
wire na1433_6;
wire na1434_1;
wire na1434_2;
wire na1434_4;
wire na1434_7;
wire na1435_1;
wire na1435_3_i;
wire na1435_4;
wire na1435_5;
wire na1435_7;
wire na1436_3;
wire na1436_4;
wire na1436_5;
wire na1436_7;
wire na1437_1;
wire na1437_2;
wire na1437_3;
wire na1437_3_i;
wire na1437_4;
wire na1437_5;
wire na1437_7;
wire na1437_8;
wire na1438_4;
wire na1438_5;
wire na1438_7;
wire na1438_8;
wire na1439_3;
wire na1439_4;
wire na1439_5;
wire na1439_6;
wire na1439_7;
wire na1439_8;
wire na1440_3;
wire na1440_4;
wire na1440_5;
wire na1440_6;
wire na1440_7;
wire na1440_8;
wire na1441_3;
wire na1441_4;
wire na1441_5;
wire na1441_6;
wire na1441_7;
wire na1441_8;
wire na1442_3;
wire na1442_4;
wire na1442_5;
wire na1442_6;
wire na1442_7;
wire na1442_8;
wire na1443_3;
wire na1443_4;
wire na1443_5;
wire na1443_6;
wire na1443_7;
wire na1443_8;
wire na1444_3;
wire na1444_4;
wire na1444_5;
wire na1444_6;
wire na1444_7;
wire na1444_8;
wire na1445_3;
wire na1445_4;
wire na1445_5;
wire na1445_6;
wire na1445_7;
wire na1445_8;
wire na1446_3;
wire na1446_4;
wire na1446_5;
wire na1446_6;
wire na1446_7;
wire na1446_8;
wire na1447_3;
wire na1447_4;
wire na1447_5;
wire na1447_6;
wire na1447_7;
wire na1447_8;
wire na1448_3;
wire na1448_4;
wire na1448_5;
wire na1448_6;
wire na1448_7;
wire na1448_8;
wire na1449_3;
wire na1449_4;
wire na1449_5;
wire na1449_6;
wire na1449_7;
wire na1449_8;
wire na1450_3;
wire na1450_4;
wire na1450_5;
wire na1450_6;
wire na1450_7;
wire na1450_8;
wire na1451_3;
wire na1451_4;
wire na1451_5;
wire na1451_6;
wire na1451_7;
wire na1451_8;
wire na1452_3;
wire na1452_4;
wire na1452_5;
wire na1452_6;
wire na1452_7;
wire na1452_8;
wire na1453_3;
wire na1453_4;
wire na1453_5;
wire na1453_6;
wire na1453_7;
wire na1453_8;
wire na1454_3;
wire na1454_4;
wire na1454_5;
wire na1454_6;
wire na1454_7;
wire na1454_8;
wire na1455_2;
wire na1455_3;
wire na1455_3_i;
wire na1455_6;
wire na1456_1;
wire na1456_2;
wire na1456_4;
wire na1456_7;
wire na1457_1;
wire na1457_3_i;
wire na1457_4;
wire na1457_5;
wire na1457_7;
wire na1458_3;
wire na1458_4;
wire na1458_5;
wire na1458_7;
wire na1459_1;
wire na1459_2;
wire na1459_3;
wire na1459_3_i;
wire na1459_4;
wire na1459_5;
wire na1459_7;
wire na1459_8;
wire na1460_4;
wire na1460_5;
wire na1460_7;
wire na1460_8;
wire na1461_3;
wire na1461_4;
wire na1461_5;
wire na1461_6;
wire na1461_7;
wire na1461_8;
wire na1462_3;
wire na1462_4;
wire na1462_5;
wire na1462_6;
wire na1462_7;
wire na1462_8;
wire na1463_3;
wire na1463_4;
wire na1463_5;
wire na1463_6;
wire na1463_7;
wire na1463_8;
wire na1464_3;
wire na1464_4;
wire na1464_5;
wire na1464_6;
wire na1464_7;
wire na1464_8;
wire na1465_3;
wire na1465_4;
wire na1465_5;
wire na1465_6;
wire na1465_7;
wire na1465_8;
wire na1466_3;
wire na1466_4;
wire na1466_5;
wire na1466_6;
wire na1466_7;
wire na1466_8;
wire na1467_3;
wire na1467_4;
wire na1467_5;
wire na1467_6;
wire na1467_7;
wire na1467_8;
wire na1468_3;
wire na1468_4;
wire na1468_5;
wire na1468_6;
wire na1468_7;
wire na1468_8;
wire na1469_3;
wire na1469_4;
wire na1469_5;
wire na1469_6;
wire na1469_7;
wire na1469_8;
wire na1470_3;
wire na1470_4;
wire na1470_5;
wire na1470_6;
wire na1470_7;
wire na1470_8;
wire na1471_3;
wire na1471_4;
wire na1471_5;
wire na1471_6;
wire na1471_7;
wire na1471_8;
wire na1472_3;
wire na1472_4;
wire na1472_5;
wire na1472_6;
wire na1472_7;
wire na1472_8;
wire na1473_3;
wire na1473_4;
wire na1473_5;
wire na1473_6;
wire na1473_7;
wire na1473_8;
wire na1474_3;
wire na1474_4;
wire na1474_5;
wire na1474_6;
wire na1474_7;
wire na1474_8;
wire na1475_3;
wire na1475_4;
wire na1475_5;
wire na1475_6;
wire na1475_7;
wire na1475_8;
wire na1476_3;
wire na1476_4;
wire na1476_5;
wire na1476_6;
wire na1476_7;
wire na1476_8;
wire na1477_2;
wire na1477_3;
wire na1477_3_i;
wire na1477_6;
wire na1478_1;
wire na1478_2;
wire na1478_4;
wire na1478_7;
wire na1479_1;
wire na1479_3_i;
wire na1479_4;
wire na1479_5;
wire na1479_7;
wire na1480_3;
wire na1480_4;
wire na1480_5;
wire na1480_7;
wire na1481_1;
wire na1481_2;
wire na1481_3;
wire na1481_3_i;
wire na1481_4;
wire na1481_5;
wire na1481_7;
wire na1481_8;
wire na1482_1;
wire na1482_2;
wire na1482_4;
wire na1482_5;
wire na1482_7;
wire na1482_8;
wire na1483_3;
wire na1483_4;
wire na1483_5;
wire na1483_6;
wire na1483_7;
wire na1483_8;
wire na1484_3;
wire na1484_4;
wire na1484_5;
wire na1484_6;
wire na1484_7;
wire na1484_8;
wire na1485_3;
wire na1485_4;
wire na1485_5;
wire na1485_6;
wire na1485_7;
wire na1485_8;
wire na1486_3;
wire na1486_4;
wire na1486_5;
wire na1486_6;
wire na1486_7;
wire na1486_8;
wire na1487_3;
wire na1487_4;
wire na1487_5;
wire na1487_6;
wire na1487_7;
wire na1487_8;
wire na1488_3;
wire na1488_4;
wire na1488_5;
wire na1488_6;
wire na1488_7;
wire na1488_8;
wire na1489_3;
wire na1489_4;
wire na1489_5;
wire na1489_6;
wire na1489_7;
wire na1489_8;
wire na1490_3;
wire na1490_4;
wire na1490_5;
wire na1490_6;
wire na1490_7;
wire na1490_8;
wire na1491_3;
wire na1491_4;
wire na1491_5;
wire na1491_6;
wire na1491_7;
wire na1491_8;
wire na1492_3;
wire na1492_4;
wire na1492_5;
wire na1492_6;
wire na1492_7;
wire na1492_8;
wire na1493_3;
wire na1493_4;
wire na1493_5;
wire na1493_6;
wire na1493_7;
wire na1493_8;
wire na1494_3;
wire na1494_4;
wire na1494_5;
wire na1494_6;
wire na1494_7;
wire na1494_8;
wire na1495_3;
wire na1495_4;
wire na1495_5;
wire na1495_6;
wire na1495_7;
wire na1495_8;
wire na1496_3;
wire na1496_4;
wire na1496_5;
wire na1496_6;
wire na1496_7;
wire na1496_8;
wire na1497_3;
wire na1497_4;
wire na1497_5;
wire na1497_6;
wire na1497_7;
wire na1497_8;
wire na1498_3;
wire na1498_4;
wire na1498_5;
wire na1498_6;
wire na1498_7;
wire na1498_8;
wire na1499_2;
wire na1499_3;
wire na1499_3_i;
wire na1499_6;
wire na1500_1;
wire na1500_2;
wire na1500_4;
wire na1500_7;
wire na1501_1;
wire na1501_3_i;
wire na1501_4;
wire na1501_5;
wire na1501_7;
wire na1502_4;
wire na1502_5;
wire na1502_7;
wire na1503_1;
wire na1503_2;
wire na1503_3_i;
wire na1503_4;
wire na1503_5;
wire na1503_7;
wire na1503_8;
wire na1504_1;
wire na1504_2;
wire na1504_4;
wire na1504_5;
wire na1504_7;
wire na1504_8;
wire na1505_1;
wire na1505_2;
wire na1505_4;
wire na1505_5;
wire na1505_7;
wire na1505_8;
wire na1506_1;
wire na1506_2;
wire na1506_4;
wire na1506_5;
wire na1506_7;
wire na1506_8;
wire na1507_1;
wire na1507_2;
wire na1507_4;
wire na1507_5;
wire na1507_7;
wire na1507_8;
wire na1508_1;
wire na1508_2;
wire na1508_4;
wire na1508_5;
wire na1508_7;
wire na1508_8;
wire na1509_1;
wire na1509_2;
wire na1509_4;
wire na1509_5;
wire na1509_7;
wire na1509_8;
wire na1510_1;
wire na1510_2;
wire na1510_4;
wire na1510_5;
wire na1510_7;
wire na1510_8;
wire na1511_1;
wire na1511_2;
wire na1511_4;
wire na1511_5;
wire na1511_7;
wire na1511_8;
wire na1512_1;
wire na1512_2;
wire na1512_4;
wire na1512_5;
wire na1512_7;
wire na1512_8;
wire na1513_1;
wire na1513_2;
wire na1513_4;
wire na1513_5;
wire na1513_7;
wire na1513_8;
wire na1514_1;
wire na1514_2;
wire na1514_4;
wire na1514_5;
wire na1514_7;
wire na1514_8;
wire na1515_1;
wire na1515_2;
wire na1515_4;
wire na1515_5;
wire na1515_7;
wire na1515_8;
wire na1516_1;
wire na1516_2;
wire na1516_4;
wire na1516_5;
wire na1516_7;
wire na1516_8;
wire na1517_4;
wire na1517_5;
wire na1517_7;
wire na1517_8;
wire na1518_4;
wire na1518_5;
wire na1518_7;
wire na1518_8;
wire na1519_4;
wire na1519_5;
wire na1519_7;
wire na1519_8;
wire na1520_4;
wire na1520_5;
wire na1520_7;
wire na1520_8;
wire na1521_3_i;
wire na1522_2;
wire na1523_1;
wire na1523_2;
wire na1523_3;
wire na1523_3_i;
wire na1523_6;
wire na1524_1;
wire na1524_2;
wire na1524_3;
wire na1524_3_i;
wire na1524_6;
wire na1525_1;
wire na1525_2;
wire na1525_3;
wire na1525_3_i;
wire na1525_6;
wire na1526_1;
wire na1526_2;
wire na1526_3;
wire na1526_3_i;
wire na1526_6;
wire na1527_1;
wire na1527_2;
wire na1527_3;
wire na1527_3_i;
wire na1527_6;
wire na1528_1;
wire na1528_2;
wire na1528_3;
wire na1528_3_i;
wire na1528_6;
wire na1529_1;
wire na1529_2;
wire na1529_3;
wire na1529_3_i;
wire na1529_6;
wire na1530_1;
wire na1530_2;
wire na1530_3;
wire na1530_3_i;
wire na1530_6;
wire na1531_1;
wire na1531_2;
wire na1531_3;
wire na1531_3_i;
wire na1531_6;
wire na1532_1;
wire na1532_2;
wire na1532_4;
wire na1532_7;
wire na1533_1;
wire na1533_3_i;
wire na1533_4;
wire na1533_5;
wire na1533_7;
wire na1534_3;
wire na1534_4;
wire na1534_5;
wire na1534_7;
wire na1535_1;
wire na1535_2;
wire na1535_3;
wire na1535_3_i;
wire na1535_4;
wire na1535_5;
wire na1535_7;
wire na1535_8;
wire na1536_4;
wire na1536_5;
wire na1536_7;
wire na1536_8;
wire na1537_3;
wire na1537_4;
wire na1537_5;
wire na1537_6;
wire na1537_7;
wire na1537_8;
wire na1538_3;
wire na1538_4;
wire na1538_5;
wire na1538_6;
wire na1538_7;
wire na1538_8;
wire na1539_3;
wire na1539_4;
wire na1539_5;
wire na1539_6;
wire na1539_7;
wire na1539_8;
wire na1540_3;
wire na1540_4;
wire na1540_5;
wire na1540_6;
wire na1540_7;
wire na1540_8;
wire na1541_3;
wire na1541_4;
wire na1541_5;
wire na1541_6;
wire na1541_7;
wire na1541_8;
wire na1542_3;
wire na1542_4;
wire na1542_5;
wire na1542_6;
wire na1542_7;
wire na1542_8;
wire na1543_3;
wire na1543_4;
wire na1543_5;
wire na1543_6;
wire na1543_7;
wire na1543_8;
wire na1544_3;
wire na1544_4;
wire na1544_5;
wire na1544_6;
wire na1544_7;
wire na1544_8;
wire na1545_2;
wire na1545_3;
wire na1545_3_i;
wire na1545_6;
wire na1546_1;
wire na1546_2;
wire na1546_4;
wire na1546_7;
wire na1547_1;
wire na1547_3_i;
wire na1547_4;
wire na1547_5;
wire na1547_7;
wire na1548_3;
wire na1548_4;
wire na1548_5;
wire na1548_7;
wire na1549_1;
wire na1549_2;
wire na1549_3;
wire na1549_3_i;
wire na1549_4;
wire na1549_5;
wire na1549_7;
wire na1549_8;
wire na1550_4;
wire na1550_5;
wire na1550_7;
wire na1550_8;
wire na1551_3;
wire na1551_4;
wire na1551_5;
wire na1551_6;
wire na1551_7;
wire na1551_8;
wire na1552_3;
wire na1552_4;
wire na1552_5;
wire na1552_6;
wire na1552_7;
wire na1552_8;
wire na1553_3;
wire na1553_4;
wire na1553_5;
wire na1553_6;
wire na1553_7;
wire na1553_8;
wire na1554_3;
wire na1554_4;
wire na1554_5;
wire na1554_6;
wire na1554_7;
wire na1554_8;
wire na1555_3;
wire na1555_4;
wire na1555_5;
wire na1555_6;
wire na1555_7;
wire na1555_8;
wire na1556_3;
wire na1556_4;
wire na1556_5;
wire na1556_6;
wire na1556_7;
wire na1556_8;
wire na1557_3;
wire na1557_4;
wire na1557_5;
wire na1557_6;
wire na1557_7;
wire na1557_8;
wire na1558_3;
wire na1558_4;
wire na1558_5;
wire na1558_6;
wire na1558_7;
wire na1558_8;
wire na1559_2;
wire na1559_3;
wire na1559_3_i;
wire na1559_6;
wire na1560_1;
wire na1560_2;
wire na1560_4;
wire na1560_7;
wire na1561_1;
wire na1561_3_i;
wire na1561_4;
wire na1561_5;
wire na1561_7;
wire na1562_3;
wire na1562_4;
wire na1562_5;
wire na1562_7;
wire na1563_1;
wire na1563_2;
wire na1563_3;
wire na1563_3_i;
wire na1563_4;
wire na1563_5;
wire na1563_7;
wire na1563_8;
wire na1564_4;
wire na1564_5;
wire na1564_7;
wire na1564_8;
wire na1565_3;
wire na1565_4;
wire na1565_5;
wire na1565_6;
wire na1565_7;
wire na1565_8;
wire na1566_3;
wire na1566_4;
wire na1566_5;
wire na1566_6;
wire na1566_7;
wire na1566_8;
wire na1567_3;
wire na1567_4;
wire na1567_5;
wire na1567_6;
wire na1567_7;
wire na1567_8;
wire na1568_3;
wire na1568_4;
wire na1568_5;
wire na1568_6;
wire na1568_7;
wire na1568_8;
wire na1569_3;
wire na1569_4;
wire na1569_5;
wire na1569_6;
wire na1569_7;
wire na1569_8;
wire na1570_3;
wire na1570_4;
wire na1570_5;
wire na1570_6;
wire na1570_7;
wire na1570_8;
wire na1571_3;
wire na1571_4;
wire na1571_5;
wire na1571_6;
wire na1571_7;
wire na1571_8;
wire na1572_3;
wire na1572_4;
wire na1572_5;
wire na1572_6;
wire na1572_7;
wire na1572_8;
wire na1573_2;
wire na1573_3;
wire na1573_3_i;
wire na1573_6;
wire na1574_1;
wire na1574_2;
wire na1574_4;
wire na1574_7;
wire na1575_1;
wire na1575_3_i;
wire na1575_4;
wire na1575_5;
wire na1575_7;
wire na1576_3;
wire na1576_4;
wire na1576_5;
wire na1576_7;
wire na1577_1;
wire na1577_2;
wire na1577_3;
wire na1577_3_i;
wire na1577_4;
wire na1577_5;
wire na1577_7;
wire na1577_8;
wire na1578_1;
wire na1578_2;
wire na1578_4;
wire na1578_5;
wire na1578_7;
wire na1578_8;
wire na1579_3;
wire na1579_4;
wire na1579_5;
wire na1579_6;
wire na1579_7;
wire na1579_8;
wire na1580_3;
wire na1580_4;
wire na1580_5;
wire na1580_6;
wire na1580_7;
wire na1580_8;
wire na1581_3;
wire na1581_4;
wire na1581_5;
wire na1581_6;
wire na1581_7;
wire na1581_8;
wire na1582_3;
wire na1582_4;
wire na1582_5;
wire na1582_6;
wire na1582_7;
wire na1582_8;
wire na1583_3;
wire na1583_4;
wire na1583_5;
wire na1583_6;
wire na1583_7;
wire na1583_8;
wire na1584_3;
wire na1584_4;
wire na1584_5;
wire na1584_6;
wire na1584_7;
wire na1584_8;
wire na1585_3;
wire na1585_4;
wire na1585_5;
wire na1585_6;
wire na1585_7;
wire na1585_8;
wire na1586_3;
wire na1586_4;
wire na1586_5;
wire na1586_6;
wire na1586_7;
wire na1586_8;
wire na1587_2;
wire na1587_3;
wire na1587_3_i;
wire na1587_6;
wire na1588_1;
wire na1588_2;
wire na1588_4;
wire na1588_7;
wire na1589_1;
wire na1589_3_i;
wire na1589_4;
wire na1589_5;
wire na1589_7;
wire na1590_4;
wire na1590_5;
wire na1590_7;
wire na1591_1;
wire na1591_2;
wire na1591_3_i;
wire na1591_4;
wire na1591_5;
wire na1591_7;
wire na1591_8;
wire na1592_1;
wire na1592_2;
wire na1592_4;
wire na1592_5;
wire na1592_7;
wire na1592_8;
wire na1593_1;
wire na1593_2;
wire na1593_4;
wire na1593_5;
wire na1593_7;
wire na1593_8;
wire na1594_1;
wire na1594_2;
wire na1594_4;
wire na1594_5;
wire na1594_7;
wire na1594_8;
wire na1595_1;
wire na1595_2;
wire na1595_4;
wire na1595_5;
wire na1595_7;
wire na1595_8;
wire na1596_1;
wire na1596_2;
wire na1596_4;
wire na1596_5;
wire na1596_7;
wire na1596_8;
wire na1597_1;
wire na1597_2;
wire na1597_4;
wire na1597_5;
wire na1597_7;
wire na1597_8;
wire na1598_1;
wire na1598_2;
wire na1598_4;
wire na1598_5;
wire na1598_7;
wire na1598_8;
wire na1599_4;
wire na1599_5;
wire na1599_7;
wire na1599_8;
wire na1600_4;
wire na1600_5;
wire na1600_7;
wire na1600_8;
wire na1601_3_i;
wire na1602_2;
wire na1603_2;
wire na1604_2;
wire na1605_2;
wire na1606_2;
wire na1607_2;
wire na1608_2;
wire na1609_2;
wire na1610_2;
wire na1611_2;
wire na1612_2;
wire na1613_2;
wire na1614_2;
wire na1615_2;
wire na1616_2;
wire na1617_2;
wire na1618_2;
wire na1619_2;
wire na1620_2;
wire na1621_2;
wire na1622_2;
wire na1623_2;
wire na1624_2;
wire na1625_2;
wire na1626_2;
wire na1627_2;
wire na1628_2;
wire na1629_2;
wire na1630_2;
wire na1631_2;
wire na1632_2;
wire na1633_2;
wire na1634_2;
wire na1635_2;
wire na1636_2;
wire na1637_2;
wire na1638_2;
wire na1639_2;
wire na1640_2;
wire na1641_2;
wire na1642_2;
wire na1643_2;
wire na1644_2;
wire na1645_2;
wire na1646_2;
wire na1647_2;
wire na1648_2;
wire na1649_2;
wire na1650_2;
wire na1651_2;
wire na1652_2;
wire na1653_2;
wire na1654_2;
wire na1655_2;
wire na1656_2;
wire na1657_2;
wire na1658_2;
wire na1659_2;
wire na1660_2;
wire na1661_2;
wire na1662_2;
wire na1663_2;
wire na1664_2;
wire na1665_2;
wire na1666_2;
wire na1667_2;
wire na1668_2;
wire na1669_2;
wire na1670_2;
wire na1671_2;
wire na1672_2;
wire na1673_2;
wire na1674_2;
wire na1675_2;
wire na1676_2;
wire na1677_2;
wire na1678_2;
wire na1679_2;
wire na1680_2;
wire na1681_2;
wire na1682_2;
wire na1683_2;
wire na1684_2;
wire na1685_2;
wire na1686_2;
wire na1687_2;
wire na1688_2;
wire na1689_2;
wire na1690_2;
wire na1691_2;
wire na1692_2;
wire na1693_2;
wire na1694_2;
wire na1695_2;
wire na1696_2;
wire na1697_2;
wire na1698_2;
wire na1699_2;
wire na1700_2;
wire na1701_2;
wire na1702_2;
wire na1703_2;
wire na1704_2;
wire na1705_2;
wire na1706_2;
wire na1707_2;
wire na1708_2;
wire na1709_2;
wire na1710_2;
wire na1711_2;
wire na1712_2;
wire na1713_2;
wire na1714_2;
wire na1715_2;
wire na1716_2;
wire na1717_2;
wire na1718_2;
wire na1719_2;
wire na1720_2;
wire na1721_2;
wire na1722_2;
wire na1723_2;
wire na1724_2;
wire na1725_2;
wire na1726_2;
wire na1727_2;
wire na1728_2;
wire na1729_2;
wire na1730_2;
wire na1731_2;
wire na1732_2;
wire na1733_2;
wire na1734_2;
wire na1735_2;
wire na1736_2;
wire na1737_2;
wire na1738_2;
wire na1739_2;
wire na1740_2;
wire na1741_2;
wire na1742_2;
wire na1743_2;
wire na1744_2;
wire na1745_2;
wire na1746_2;
wire na1747_2;
wire na1748_2;
wire na1749_2;
wire na1750_2;
wire na1751_2;
wire na1752_2;
wire na1753_2;
wire na1754_2;
wire na1755_2;
wire na1756_2;
wire na1757_2;
wire na1758_2;
wire na1759_2;
wire na1760_2;
wire na1761_2;
wire na1762_2;
wire na1763_2;
wire na1764_2;
wire na1765_2;
wire na1766_2;
wire na1767_2;
wire na1768_2;
wire na1769_2;
wire na1770_2;
wire na1771_2;
wire na1772_2;
wire na1773_2;
wire na1774_2;
wire na1775_2;
wire na1776_2;
wire na1777_2;
wire na1778_2;
wire na1779_2;
wire na1780_2;
wire na1781_2;
wire na1782_2;
wire na1783_2;
wire na1784_2;
wire na1785_2;
wire na1786_2;
wire na1787_2;
wire na1788_2;
wire na1789_2;
wire na1790_2;
wire na1791_2;
wire na1792_2;
wire na1793_2;
wire na1794_2;
wire na1795_2;
wire na1796_2;
wire na1797_2;
wire na1798_2;
wire na1799_2;
wire na1800_2;
wire na1801_2;
wire na1802_2;
wire na1803_2;
wire na1804_2;
wire na1805_2;
wire na1806_2;
wire na1807_2;
wire na1808_2;
wire na1809_2;
wire na1810_2;
wire na1811_2;
wire na1812_2;
wire na1813_2;
wire na1814_2;
wire clk_10mhz;
wire na1602_10;
wire na1603_10;
wire na1604_10;
wire ant_433mhz;
wire wifi_gpio0;

// C_XOR////      x28y77     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a4_1 ( .OUT(na4_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na98_2), .IN7(1'b0), .IN8(na99_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x24y73     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a5_4 ( .OUT(na5_2), .IN1(1'b1), .IN2(~na98_2), .IN3(1'b1), .IN4(na99_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x21y73     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a6_1 ( .OUT(na6_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na98_2), .IN7(1'b1), .IN8(~na99_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x27y78     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a7_4 ( .OUT(na7_2), .IN1(1'b1), .IN2(na98_2), .IN3(1'b1), .IN4(~na99_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x22y79     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a8_1 ( .OUT(na8_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na98_2), .IN7(1'b1), .IN8(na99_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x23y78     80'h00_0018_00_0040_0C8E_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a9_1 ( .OUT(na9_1), .IN1(1'b0), .IN2(na1042_1), .IN3(na1799_2), .IN4(~na99_1), .IN5(1'b1), .IN6(na98_1), .IN7(1'b1), .IN8(na99_2),
                   .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x26y82     80'h00_0018_00_0040_0C09_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a10_1 ( .OUT(na10_1), .IN1(na1043_2), .IN2(1'b0), .IN3(1'b0), .IN4(na1044_1), .IN5(na1645_2), .IN6(1'b1), .IN7(1'b1), .IN8(na99_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x24y80     80'h00_0018_00_0040_0C06_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a11_1 ( .OUT(na11_1), .IN1(1'b0), .IN2(na98_1), .IN3(na1045_2), .IN4(1'b0), .IN5(1'b1), .IN6(na98_2), .IN7(1'b1), .IN8(na99_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x28y78     80'h00_0018_00_0040_0C29_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a12_1 ( .OUT(na12_1), .IN1(na1046_1), .IN2(1'b1), .IN3(1'b0), .IN4(na1047_2), .IN5(1'b1), .IN6(na98_2), .IN7(na1640_2),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x30y79     80'h00_0018_00_0040_0CEE_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a13_1 ( .OUT(na13_1), .IN1(1'b0), .IN2(~na98_1), .IN3(~na1049_2), .IN4(~na1048_1), .IN5(1'b1), .IN6(~na98_2), .IN7(1'b1),
                    .IN8(na99_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x21y75     80'h00_0018_00_0040_0AB7_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a14_1 ( .OUT(na14_1), .IN1(1'b1), .IN2(na98_1), .IN3(1'b1), .IN4(na99_2), .IN5(~na1643_2), .IN6(~na1042_1), .IN7(1'b1),
                    .IN8(na99_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x25y77     80'h00_0018_00_0040_0C1D_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a15_1 ( .OUT(na15_1), .IN1(~na6_1), .IN2(1'b0), .IN3(na1611_2), .IN4(na1606_2), .IN5(1'b1), .IN6(~na98_1), .IN7(1'b1), .IN8(~na99_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x25y80     80'h00_0018_00_0040_0AB8_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a16_1 ( .OUT(na16_1), .IN1(1'b1), .IN2(na98_1), .IN3(1'b1), .IN4(na99_2), .IN5(na1041_2), .IN6(na1054_1), .IN7(1'b0), .IN8(~na99_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x24y75     80'h00_0018_00_0040_0C92_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a17_1 ( .OUT(na17_1), .IN1(1'b1), .IN2(na7_2), .IN3(1'b0), .IN4(1'b1), .IN5(1'b1), .IN6(~na98_1), .IN7(1'b1), .IN8(na99_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x31y77     80'h00_0018_00_0040_0C0F_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a18_1 ( .OUT(na18_1), .IN1(na1055_2), .IN2(na98_1), .IN3(na1644_2), .IN4(na1800_2), .IN5(1'b1), .IN6(na98_2), .IN7(1'b1),
                    .IN8(~na99_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x30y80     80'h00_0060_00_0000_0C0E_FF0B
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a19_4 ( .OUT(na19_2), .IN1(na1056_1), .IN2(~na98_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x29y76     80'h00_0060_00_0000_0C08_FFF2
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a20_4 ( .OUT(na20_2), .IN1(na611_1), .IN2(~na871_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x32y73     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a21_4 ( .OUT(na21_2), .IN1(~na611_1), .IN2(na871_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x32y80     80'h00_0018_00_0000_0C66_0900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a22_1 ( .OUT(na22_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na611_1), .IN6(na871_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x52y48     80'h00_0060_00_0000_0C06_FF3C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a23_4 ( .OUT(na23_2), .IN1(1'b0), .IN2(na583_1), .IN3(1'b0), .IN4(~na866_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x48y54     80'h00_0078_00_0000_0C88_C34F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a24_1 ( .OUT(na24_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na583_1), .IN7(1'b1), .IN8(na866_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a24_4 ( .OUT(na24_2), .IN1(1'b1), .IN2(1'b1), .IN3(~na868_1), .IN4(na90_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x47y54     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a25_1 ( .OUT(na25_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na583_1), .IN7(1'b1), .IN8(na866_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x50y51     80'h00_0060_00_0000_0C08_FF33
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a26_4 ( .OUT(na26_2), .IN1(1'b1), .IN2(~na583_1), .IN3(1'b1), .IN4(~na866_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y46     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a27_1 ( .OUT(na27_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na583_1), .IN7(1'b1), .IN8(~na866_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x48y50     80'h00_0018_00_0040_0C68_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a28_1 ( .OUT(na28_1), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(na866_1), .IN5(1'b1), .IN6(na583_1), .IN7(1'b1), .IN8(na866_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x47y51     80'h00_0060_00_0000_0C06_FF60
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a29_4 ( .OUT(na29_2), .IN1(1'b0), .IN2(1'b0), .IN3(na26_2), .IN4(na866_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x48y52     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a30_1 ( .OUT(na30_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na26_2), .IN8(na866_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x49y53     80'h00_0060_00_0000_0C08_FF35
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a31_4 ( .OUT(na31_2), .IN1(~na1739_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na27_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND///ORAND/      x50y47     80'h00_0078_00_0000_0C88_37CE
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a32_1 ( .OUT(na32_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1739_2), .IN6(~na583_1), .IN7(1'b0), .IN8(~na866_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a32_4 ( .OUT(na32_2), .IN1(na585_1), .IN2(na1742_2), .IN3(1'b0), .IN4(na90_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x36y68     80'h00_FA00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a35_1 ( .OUT(na35_1_i), .IN1(1'b1), .IN2(~na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na444_1), .IN6(na1681_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a35_2 ( .OUT(na35_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na35_1_i) );
// C_MX2b/D///      x33y69     80'h00_FA00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a36_1 ( .OUT(na36_1_i), .IN1(1'b1), .IN2(~na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na444_2), .IN6(na1682_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a36_2 ( .OUT(na36_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na36_1_i) );
// C_MX2b/D///      x35y71     80'h00_FA00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a37_1 ( .OUT(na37_1_i), .IN1(1'b1), .IN2(na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1683_2), .IN6(na446_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a37_2 ( .OUT(na37_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na37_1_i) );
// C_MX2b/D///      x29y65     80'h00_FA00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a38_1 ( .OUT(na38_1_i), .IN1(1'b1), .IN2(na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1684_2), .IN6(na446_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a38_2 ( .OUT(na38_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na38_1_i) );
// C_MX2b/D///      x38y70     80'h00_FA00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a39_1 ( .OUT(na39_1_i), .IN1(1'b1), .IN2(~na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na448_1), .IN6(na1685_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a39_2 ( .OUT(na39_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na39_1_i) );
// C_MX2b/D///      x41y73     80'h00_FA00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a40_1 ( .OUT(na40_1_i), .IN1(1'b1), .IN2(~na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na448_2), .IN6(na1686_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a40_2 ( .OUT(na40_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na40_1_i) );
// C_MX2b/D///      x33y66     80'h00_FA00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a41_1 ( .OUT(na41_1_i), .IN1(1'b1), .IN2(na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1687_2), .IN6(na450_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a41_2 ( .OUT(na41_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na41_1_i) );
// C_MX2b/D///      x34y68     80'h00_FA00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a42_1 ( .OUT(na42_1_i), .IN1(1'b1), .IN2(na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1688_2), .IN6(na450_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a42_2 ( .OUT(na42_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na42_1_i) );
// C_MX2b/D///      x34y69     80'h00_FA00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a43_1 ( .OUT(na43_1_i), .IN1(1'b1), .IN2(~na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na452_1), .IN6(na1689_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a43_2 ( .OUT(na43_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na43_1_i) );
// C_MX2b/D///      x37y69     80'h00_FA00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a44_1 ( .OUT(na44_1_i), .IN1(1'b1), .IN2(~na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na452_2), .IN6(na1690_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a44_2 ( .OUT(na44_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na44_1_i) );
// C_MX2b/D///      x37y73     80'h00_FA00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a45_1 ( .OUT(na45_1_i), .IN1(1'b1), .IN2(na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1676_2), .IN6(na439_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a45_2 ( .OUT(na45_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na45_1_i) );
// C_MX2a/D///      x38y71     80'h00_FA00_00_0040_0C03_0C00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a46_1 ( .OUT(na46_1_i), .IN1(na1677_2), .IN2(na439_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na948_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a46_2 ( .OUT(na46_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na46_1_i) );
// C_MX2b/D///      x37y75     80'h00_FA00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a47_1 ( .OUT(na47_1_i), .IN1(1'b1), .IN2(~na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na441_1), .IN6(na1678_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a47_2 ( .OUT(na47_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na47_1_i) );
// C_MX2b/D///      x36y73     80'h00_FA00_00_0040_0A30_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a48_1 ( .OUT(na48_1_i), .IN1(1'b1), .IN2(~na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na441_2), .IN6(na1679_2), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a48_2 ( .OUT(na48_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na48_1_i) );
// C_MX2b/D///      x31y73     80'h00_FA00_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a49_1 ( .OUT(na49_1_i), .IN1(1'b1), .IN2(na948_1), .IN3(1'b0), .IN4(1'b0), .IN5(na1680_2), .IN6(na443_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a49_2 ( .OUT(na49_1), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na49_1_i) );
// C_AND///AND/      x50y53     80'h00_0078_00_0000_0C88_3A8F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a50_1 ( .OUT(na50_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1739_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na24_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a50_4 ( .OUT(na50_2), .IN1(1'b1), .IN2(1'b1), .IN3(na868_1), .IN4(na90_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x51y52     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a51_1 ( .OUT(na51_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na583_1), .IN7(1'b1), .IN8(~na866_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x54y50     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a52_4 ( .OUT(na52_2), .IN1(1'b1), .IN2(~na51_1), .IN3(1'b1), .IN4(na866_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x49y46     80'h00_0018_00_0040_0CBD_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a53_1 ( .OUT(na53_1), .IN1(~na1739_2), .IN2(1'b1), .IN3(na1741_2), .IN4(~na866_1), .IN5(1'b1), .IN6(~na583_1), .IN7(1'b1),
                    .IN8(na866_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x50y49     80'h00_0018_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a54_1 ( .OUT(na54_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na51_1), .IN7(na32_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x53y50     80'h00_0018_00_0040_0C79_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a55_1 ( .OUT(na55_1), .IN1(~na1739_2), .IN2(1'b1), .IN3(1'b1), .IN4(na866_1), .IN5(~na585_1), .IN6(1'b1), .IN7(na26_2),
                    .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x44y51     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a56_1 ( .OUT(na56_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na25_1), .IN7(1'b1), .IN8(~na866_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y75     80'h00_0018_00_0000_0C88_F1FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a57_1 ( .OUT(na57_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na611_1), .IN6(~na871_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x32y80     80'h00_0060_00_0000_0C08_FFF8
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a58_4 ( .OUT(na58_2), .IN1(na611_1), .IN2(na871_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x34y76     80'h00_0018_00_0040_0C92_3500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a60_1 ( .OUT(na60_1), .IN1(1'b1), .IN2(na871_1), .IN3(1'b0), .IN4(1'b1), .IN5(~na611_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1746_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x36y75     80'h00_0018_00_0040_0A31_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a61_1 ( .OUT(na61_1), .IN1(1'b1), .IN2(~na613_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na62_1), .IN6(na576_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y73     80'h00_0018_00_0000_0C88_3CFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a62_1 ( .OUT(na62_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na871_2), .IN7(1'b1), .IN8(~na58_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x44y76     80'h00_0018_00_0040_0C03_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a63_1 ( .OUT(na63_1), .IN1(na64_2), .IN2(na576_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na613_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x29y77     80'h00_0060_00_0000_0C08_FFA9
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a64_4 ( .OUT(na64_2), .IN1(na1745_2), .IN2(na871_1), .IN3(~na1701_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x36y77     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a65_1 ( .OUT(na65_1), .IN1(1'b1), .IN2(na613_1), .IN3(1'b0), .IN4(1'b0), .IN5(na578_1), .IN6(~na66_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x31y78     80'h00_0018_00_0040_0C91_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a66_1 ( .OUT(na66_1), .IN1(~na611_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b1), .IN5(1'b1), .IN6(na871_1), .IN7(1'b1), .IN8(~na1746_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x37y79     80'h00_0018_00_0040_0A30_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a67_1 ( .OUT(na67_1), .IN1(1'b1), .IN2(na613_1), .IN3(1'b0), .IN4(1'b0), .IN5(na578_2), .IN6(na68_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x27y78     80'h00_0018_00_0000_0C88_39FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a68_1 ( .OUT(na68_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na611_1), .IN6(~na871_2), .IN7(1'b0), .IN8(na1744_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x38y77     80'h00_0018_00_0040_0C13_0300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a69_1 ( .OUT(na69_1), .IN1(~na70_1), .IN2(na580_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na613_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x31y79     80'h00_0018_00_0040_0CB2_3A00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a70_1 ( .OUT(na70_1), .IN1(1'b1), .IN2(~na871_1), .IN3(1'b0), .IN4(1'b1), .IN5(na611_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1746_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/D      x54y53     80'h00_FD00_80_0000_0C06_FF53
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a72_4 ( .OUT(na72_2_i), .IN1(1'b0), .IN2(~na82_1), .IN3(~na590_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a72_5 ( .OUT(na72_2), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na72_2_i) );
// C_MX2b/D///      x55y53     80'h00_FD00_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a73_1 ( .OUT(na73_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1638_2), .IN5(na601_1), .IN6(1'b0), .IN7(na590_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a73_2 ( .OUT(na73_1), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na73_1_i) );
// C_MX2a/D///      x53y56     80'h00_FD00_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a74_1 ( .OUT(na74_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1694_2), .IN4(na592_1), .IN5(1'b1), .IN6(~na82_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a74_2 ( .OUT(na74_1), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na74_1_i) );
// C_MX2b/D///      x54y54     80'h00_FD00_00_0040_0AA0_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a75_1 ( .OUT(na75_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na1638_2), .IN5(1'b0), .IN6(na603_1), .IN7(1'b0), .IN8(na592_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a75_2 ( .OUT(na75_1), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na75_1_i) );
// C_MX2b/D///      x54y56     80'h00_FD00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a76_1 ( .OUT(na76_1_i), .IN1(1'b1), .IN2(na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na594_1), .IN8(na1695_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a76_2 ( .OUT(na76_1), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na76_1_i) );
// C_MX2b/D///      x54y58     80'h00_FD00_00_0040_0A50_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a77_1 ( .OUT(na77_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1638_2), .IN5(na605_1), .IN6(1'b0), .IN7(na594_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a77_2 ( .OUT(na77_1), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na77_1_i) );
// C_MX2b/D///      x48y55     80'h00_FD00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a78_1 ( .OUT(na78_1_i), .IN1(1'b1), .IN2(~na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1696_2), .IN8(na596_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a78_2 ( .OUT(na78_1), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na78_1_i) );
// C_MX2a/D///      x57y58     80'h00_FD00_00_0040_0C0C_F300
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a79_1 ( .OUT(na79_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na1697_2), .IN4(na596_2), .IN5(1'b1), .IN6(~na82_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a79_2 ( .OUT(na79_1), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na79_1_i) );
// C_MX2b/D///      x53y64     80'h00_FD00_00_0040_0AC0_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a80_1 ( .OUT(na80_1_i), .IN1(1'b1), .IN2(na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na598_1), .IN8(na1698_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a80_2 ( .OUT(na80_1), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na80_1_i) );
// C_MX2a/D///      x54y60     80'h00_FD00_00_0040_0C0C_FC00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a81_1 ( .OUT(na81_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(na598_2), .IN4(na1699_2), .IN5(1'b1), .IN6(na82_1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a81_2 ( .OUT(na81_1), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na81_1_i) );
// C_MX2b/D///      x45y56     80'h00_FD00_00_0040_0AC0_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a82_1 ( .OUT(na82_1_i), .IN1(1'b1), .IN2(~na82_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na1700_2), .IN8(na589_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a82_2 ( .OUT(na82_1), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na82_1_i) );
// C_MX2b/D///      x28y73     80'h00_FA00_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a83_1 ( .OUT(na83_1_i), .IN1(na84_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na93_1), .IN6(na993_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a83_2 ( .OUT(na83_1), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na83_1_i) );
// C_///AND/      x29y69     80'h00_0060_00_0000_0C08_FF8C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a84_4 ( .OUT(na84_2), .IN1(1'b1), .IN2(na1738_2), .IN3(na426_1), .IN4(na862_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b/D///      x21y72     80'h00_FA00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a85_1 ( .OUT(na85_1_i), .IN1(na84_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na83_1), .IN8(na996_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a85_2 ( .OUT(na85_1), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na85_1_i) );
// C_MX2b/D///      x27y71     80'h00_FA00_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a86_1 ( .OUT(na86_1_i), .IN1(~na84_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na998_1), .IN6(na85_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a86_2 ( .OUT(na86_1), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na86_1_i) );
// C_MX2b/D///      x29y74     80'h00_FA00_00_0040_0A30_000A
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a87_1 ( .OUT(na87_1_i), .IN1(na84_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na86_1), .IN6(na1001_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a87_2 ( .OUT(na87_1), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na87_1_i) );
// C_MX2b/D///      x27y72     80'h00_FA00_00_0040_0A30_0005
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a88_1 ( .OUT(na88_1_i), .IN1(~na84_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na1004_1), .IN6(na87_1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a88_2 ( .OUT(na88_1), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na88_1_i) );
// C_MX2a/D///      x32y69     80'h00_FA00_00_0040_0C03_0500
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a89_1 ( .OUT(na89_1_i), .IN1(na1007_1), .IN2(na88_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na84_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a89_2 ( .OUT(na89_1), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na89_1_i) );
// C_MX2b/D///      x46y62     80'h00_FA00_00_0040_0AC0_00FA
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a90_1 ( .OUT(na90_1_i), .IN1(na84_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(na89_1), .IN8(na1009_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a90_2 ( .OUT(na90_1), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na90_1_i) );
// C_XOR/D//AND/D      x33y73     80'h00_FA00_80_0000_0C68_A55A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a91_1 ( .OUT(na91_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na91_1), .IN6(1'b0), .IN7(na1639_2), .IN8(1'b0),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a91_2 ( .OUT(na91_1), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na91_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a91_4 ( .OUT(na91_2_i), .IN1(na91_1), .IN2(1'b1), .IN3(~na1639_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a91_5 ( .OUT(na91_2), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na91_2_i) );
// C_AND/D///      x25y73     80'h00_FA00_00_0000_0C88_AAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a93_1 ( .OUT(na93_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na84_2), .IN6(1'b1), .IN7(na990_1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a93_2 ( .OUT(na93_1), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na93_1_i) );
// C_///AND/D      x20y76     80'h00_FA00_80_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a94_4 ( .OUT(na94_2_i), .IN1(~na95_1), .IN2(1'b1), .IN3(na545_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a94_5 ( .OUT(na94_2), .CLK(na624_1), .EN(na167_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na94_2_i) );
// C_AND////      x25y79     80'h00_0018_00_0000_0888_CA23
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a95_1 ( .OUT(na95_1), .IN1(1'b1), .IN2(~na98_1), .IN3(na8_1), .IN4(~na99_1), .IN5(na97_1), .IN6(1'b1), .IN7(1'b1), .IN8(na94_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND/D///      x23y75     80'h00_FA00_00_0000_0C88_C5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a97_1 ( .OUT(na97_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na95_1), .IN6(1'b1), .IN7(1'b1), .IN8(na543_2),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a97_2 ( .OUT(na97_1), .CLK(na624_1), .EN(na167_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na97_1_i) );
// C_AND/D//AND/D      x23y80     80'h00_FA00_80_0000_0C88_C5A5
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a98_1 ( .OUT(na98_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na95_1), .IN6(1'b1), .IN7(1'b1), .IN8(na543_1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a98_2 ( .OUT(na98_1), .CLK(na624_1), .EN(na167_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na98_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a98_4 ( .OUT(na98_2_i), .IN1(~na95_1), .IN2(1'b1), .IN3(na541_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a98_5 ( .OUT(na98_2), .CLK(na624_1), .EN(na167_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na98_2_i) );
// C_AND/D//AND/D      x30y78     80'h00_FA00_80_0000_0C88_A535
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a99_1 ( .OUT(na99_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na95_1), .IN6(1'b1), .IN7(na541_2), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a99_2 ( .OUT(na99_1), .CLK(na624_1), .EN(na167_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na99_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a99_4 ( .OUT(na99_2_i), .IN1(~na95_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na99_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                    .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a99_5 ( .OUT(na99_2), .CLK(na624_1), .EN(na167_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na99_2_i) );
// C_AND////      x25y53     80'h00_0018_00_0000_0888_1351
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a103_1 ( .OUT(na103_1), .IN1(~na106_2), .IN2(~na109_1), .IN3(~na110_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na109_2), .IN7(~na110_1),
                     .IN8(~na107_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND*/D      x25y55     80'h00_FA00_80_0000_0C07_FF55
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a106_4 ( .OUT(na106_2_i), .IN1(~na103_1), .IN2(1'b1), .IN3(~na549_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a106_5 ( .OUT(na106_2), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na106_2_i) );
// C_AND*/D///      x24y52     80'h00_FA00_00_0000_0388_35FF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a107_1 ( .OUT(na107_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na103_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na547_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a107_2 ( .OUT(na107_1), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na107_1_i) );
// C_///AND/D      x52y73     80'h00_FA00_80_0000_0C08_FFCA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a108_4 ( .OUT(na108_2_i), .IN1(na502_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1032_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a108_5 ( .OUT(na108_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na108_2_i) );
// C_AND*/D//AND/D      x25y56     80'h00_FA00_80_0000_0388_F4A5
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a109_1 ( .OUT(na109_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na103_1), .IN6(na109_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a109_2 ( .OUT(na109_1), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na109_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a109_4 ( .OUT(na109_2_i), .IN1(~na103_1), .IN2(1'b1), .IN3(na549_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a109_5 ( .OUT(na109_2), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na109_2_i) );
// C_AND*/D//AND*/D      x22y53     80'h00_FA00_80_0000_0387_3535
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a110_1 ( .OUT(na110_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na103_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na547_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a110_2 ( .OUT(na110_1), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na110_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a110_4 ( .OUT(na110_2_i), .IN1(~na103_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na551_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a110_5 ( .OUT(na110_2), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na110_2_i) );
// C_AND/D///      x60y69     80'h00_FA00_00_0000_0C88_8FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a111_1 ( .OUT(na111_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na704_2), .IN8(na1032_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a111_2 ( .OUT(na111_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na111_1_i) );
// C_AND/D///      x52y67     80'h00_FA00_00_0000_0C88_CAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a112_1 ( .OUT(na112_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na498_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1032_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a112_2 ( .OUT(na112_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na112_1_i) );
// C_///AND/D      x56y72     80'h00_FA00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a113_4 ( .OUT(na113_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na706_1), .IN4(na1032_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a113_5 ( .OUT(na113_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na113_2_i) );
// C_AND/D///      x50y72     80'h00_FA00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a114_1 ( .OUT(na114_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na500_1), .IN7(1'b1), .IN8(na1032_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a114_2 ( .OUT(na114_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na114_1_i) );
// C_///AND/D      x56y71     80'h00_FA00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a115_4 ( .OUT(na115_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1032_1), .IN4(na708_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a115_5 ( .OUT(na115_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na115_2_i) );
// C_AND/D//AND/D      x52y72     80'h00_FA00_80_0000_0C88_CACA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a116_1 ( .OUT(na116_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na509_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1032_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a116_2 ( .OUT(na116_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na116_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a116_4 ( .OUT(na116_2_i), .IN1(na1032_1), .IN2(1'b1), .IN3(1'b1), .IN4(na702_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a116_5 ( .OUT(na116_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na116_2_i) );
// C_AND/D///      x55y67     80'h00_FA00_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a118_1 ( .OUT(na118_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na511_1), .IN7(1'b1), .IN8(na1032_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a118_2 ( .OUT(na118_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na118_1_i) );
// C_///AND/D      x56y69     80'h00_FA00_80_0000_0C08_FF8F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a119_4 ( .OUT(na119_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na1032_1), .IN4(na700_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a119_5 ( .OUT(na119_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na119_2_i) );
// C_XOR////      x55y71     80'h00_0018_00_0000_0C66_C900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a120_1 ( .OUT(na120_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1647_2), .IN6(na889_1), .IN7(1'b0), .IN8(na121_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x56y68     80'h00_0018_00_0040_0C29_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a121_1 ( .OUT(na121_1), .IN1(na1777_2), .IN2(1'b1), .IN3(1'b0), .IN4(na967_1), .IN5(~na1650_2), .IN6(1'b1), .IN7(1'b1), .IN8(na957_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x57y69     80'h00_0018_00_0000_0666_A55E
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a122_1 ( .OUT(na122_1), .IN1(~na1647_2), .IN2(~na889_1), .IN3(na965_1), .IN4(1'b1), .IN5(na1648_2), .IN6(1'b1), .IN7(~na969_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x53y67     80'h00_0060_00_0000_0C06_FF69
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a124_4 ( .OUT(na124_2), .IN1(~na118_1), .IN2(na891_1), .IN3(na1749_2), .IN4(na1060_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x45y72     80'h00_0060_00_0000_0C06_FFA9
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a125_4 ( .OUT(na125_2), .IN1(~na118_1), .IN2(na891_1), .IN3(na1749_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x56y71     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a127_1 ( .OUT(na127_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1781_2), .IN7(~na111_1), .IN8(na967_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x56y74     80'h00_0078_00_0000_0C66_9696
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a128_1 ( .OUT(na128_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1062_1), .IN6(na893_1), .IN7(~na112_1), .IN8(na1752_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a128_4 ( .OUT(na128_2), .IN1(na1061_1), .IN2(na1781_2), .IN3(~na111_1), .IN4(na967_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x60y74     80'h00_0060_00_0000_0C06_FF56
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a129_4 ( .OUT(na129_2), .IN1(na897_1), .IN2(na893_1), .IN3(~na112_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x56y73     80'h00_0018_00_0000_0C66_9A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a131_1 ( .OUT(na131_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1769_2), .IN6(1'b0), .IN7(na969_1), .IN8(~na113_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x55y73     80'h00_0078_00_0000_0C66_9696
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a132_1 ( .OUT(na132_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1064_1), .IN6(na899_1), .IN7(na1749_2), .IN8(~na114_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a132_4 ( .OUT(na132_2), .IN1(na1769_2), .IN2(na1063_1), .IN3(na969_1), .IN4(~na113_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x50y71     80'h00_0060_00_0000_0C06_FF36
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a133_4 ( .OUT(na133_2), .IN1(na895_1), .IN2(na899_1), .IN3(1'b0), .IN4(~na114_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x55y74     80'h00_0018_00_0000_0C66_9A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a135_1 ( .OUT(na135_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1771_2), .IN6(1'b0), .IN7(~na115_2), .IN8(na971_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x55y72     80'h00_0078_00_0000_0C66_9696
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a136_1 ( .OUT(na136_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1066_1), .IN6(na901_1), .IN7(~na108_2), .IN8(na1752_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a136_4 ( .OUT(na136_2), .IN1(na1065_1), .IN2(na1772_2), .IN3(~na115_2), .IN4(na971_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x44y80     80'h00_0060_00_0000_0C06_FF56
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a137_4 ( .OUT(na137_2), .IN1(na897_1), .IN2(na901_1), .IN3(~na108_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x49y64     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a138_1 ( .OUT(na138_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na139_1), .IN7(na721_2), .IN8(~na116_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x59y70     80'h00_0018_00_0040_0C16_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a139_1 ( .OUT(na139_1), .IN1(1'b1), .IN2(na983_1), .IN3(na1792_2), .IN4(1'b0), .IN5(1'b1), .IN6(na973_1), .IN7(na119_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x59y71     80'h00_0018_00_0000_0666_3AE5
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a140_1 ( .OUT(na140_1), .IN1(na981_1), .IN2(1'b1), .IN3(~na721_2), .IN4(~na116_1), .IN5(~na985_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na116_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x54y68     80'h00_0018_00_0000_0C66_6900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a142_1 ( .OUT(na142_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na118_1), .IN6(na727_2), .IN7(na1067_1), .IN8(na723_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x60y72     80'h00_0018_00_0000_0C66_C900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a143_1 ( .OUT(na143_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na118_1), .IN6(na727_2), .IN7(1'b0), .IN8(na723_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x57y70     80'h00_0060_00_0000_0C06_FF9C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a145_4 ( .OUT(na145_2), .IN1(1'b0), .IN2(na983_1), .IN3(~na111_1), .IN4(na1796_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x55y65     80'h00_0078_00_0000_0C66_9696
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a146_1 ( .OUT(na146_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1069_1), .IN6(na729_2), .IN7(~na112_1), .IN8(na725_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a146_4 ( .OUT(na146_2), .IN1(na1068_1), .IN2(na983_1), .IN3(~na111_1), .IN4(na1798_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x50y73     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a147_1 ( .OUT(na147_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na729_2), .IN7(~na112_1), .IN8(na725_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x55y71     80'h00_0060_00_0000_0C06_FF9A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a149_4 ( .OUT(na149_2), .IN1(na985_1), .IN2(1'b0), .IN3(na1783_2), .IN4(~na113_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x52y76     80'h00_0078_00_0000_0C66_9696
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a150_1 ( .OUT(na150_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1071_1), .IN6(na727_2), .IN7(na731_2), .IN8(~na114_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a150_4 ( .OUT(na150_2), .IN1(na985_1), .IN2(na1070_1), .IN3(na1783_2), .IN4(~na113_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x49y70     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a151_1 ( .OUT(na151_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na727_2), .IN7(na731_2), .IN8(~na114_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x56y77     80'h00_0060_00_0000_0C06_FF9C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a153_4 ( .OUT(na153_2), .IN1(1'b0), .IN2(na987_1), .IN3(~na115_2), .IN4(na1787_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x57y73     80'h00_0078_00_0000_0C66_9696
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a154_1 ( .OUT(na154_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1073_1), .IN6(na729_2), .IN7(~na108_2), .IN8(na733_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a154_4 ( .OUT(na154_2), .IN1(na1785_2), .IN2(na987_1), .IN3(~na115_2), .IN4(na1072_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x52y75     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a155_1 ( .OUT(na155_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na729_2), .IN7(~na108_2), .IN8(na733_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x35y67     80'h00_0018_00_0000_0888_5C13
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a156_1 ( .OUT(na156_1), .IN1(1'b1), .IN2(~na1675_2), .IN3(~na157_1), .IN4(~na436_1), .IN5(1'b1), .IN6(na745_2), .IN7(~na434_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x46y61     80'h00_0018_00_0000_0888_4181
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a157_1 ( .OUT(na157_1), .IN1(~na951_1), .IN2(~na948_1), .IN3(na162_2), .IN4(na161_1), .IN5(~na951_2), .IN6(~na953_2), .IN7(~na1767_2),
                     .IN8(na161_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x48y62     80'h00_0078_00_0000_0C88_1111
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a161_1 ( .OUT(na161_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na944_2), .IN6(~na946_1), .IN7(~na1764_2),
                     .IN8(~na1763_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a161_4 ( .OUT(na161_2), .IN1(~na251_1), .IN2(~na949_2), .IN3(~na1765_2), .IN4(~na173_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x48y61     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a162_4 ( .OUT(na162_2), .IN1(~na955_2), .IN2(~na942_2), .IN3(~na1762_2), .IN4(~na1768_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x48y56     80'h00_0018_00_0040_0CAA_4F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a164_1 ( .OUT(na164_1), .IN1(1'b0), .IN2(~na1010_1), .IN3(1'b0), .IN4(~na1011_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na868_1),
                     .IN8(na90_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2a////      x47y53     80'h00_0018_00_0040_0CAA_4F00
C_MX2a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a165_1 ( .OUT(na165_1), .IN1(1'b0), .IN2(~na1012_1), .IN3(1'b0), .IN4(~na1013_1), .IN5(1'b1), .IN6(1'b1), .IN7(~na868_1),
                     .IN8(na90_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR/D///      x45y54     80'h00_FA00_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a166_1 ( .OUT(na166_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na166_1), .IN7(1'b0), .IN8(na90_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a166_2 ( .OUT(na166_1), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na166_1_i) );
// C_AND////      x23y72     80'h00_0018_00_0000_0C88_12FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a167_1 ( .OUT(na167_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na168_1), .IN6(~na1738_2), .IN7(~na426_1), .IN8(~na862_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x33y65     80'h00_0018_00_0000_0888_8CF8
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a168_1 ( .OUT(na168_1), .IN1(na585_1), .IN2(na169_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na25_1), .IN7(na868_1), .IN8(na866_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x43y52     80'h00_0018_00_0000_0C88_F8FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a169_1 ( .OUT(na169_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na103_1), .IN6(na82_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x44y73     80'h00_0060_00_0000_0C08_FF54
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a171_4 ( .OUT(na171_2), .IN1(~na91_1), .IN2(na82_1), .IN3(~na1639_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x56y66     80'h00_0060_00_0000_0C08_FFAA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a172_4 ( .OUT(na172_2), .IN1(na57_1), .IN2(1'b1), .IN3(na171_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x46y64     80'h00_FE18_00_0000_0666_3506
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a173_1 ( .OUT(na173_1), .IN1(na720_1), .IN2(na844_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na1578_1), .IN6(1'b0), .IN7(1'b0), .IN8(~na925_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a173_5 ( .OUT(na173_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na173_1) );
// C_XOR///XOR/      x44y72     80'h00_0078_00_0000_0C66_C99A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a176_1 ( .OUT(na176_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1578_2), .IN6(na889_2), .IN7(1'b0), .IN8(na35_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a176_4 ( .OUT(na176_2), .IN1(na36_1), .IN2(1'b0), .IN3(na927_2), .IN4(~na1592_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y65     80'h00_0018_00_0040_0A92_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a177_1 ( .OUT(na177_1), .IN1(~na720_1), .IN2(1'b1), .IN3(1'b1), .IN4(na925_2), .IN5(na1802_2), .IN6(1'b1), .IN7(1'b0), .IN8(na1076_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x48y66     80'h00_0018_00_0040_0C29_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a178_1 ( .OUT(na178_1), .IN1(na186_1), .IN2(1'b1), .IN3(1'b0), .IN4(na1654_2), .IN5(~na1656_2), .IN6(1'b1), .IN7(na179_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y69     80'h00_0018_00_0040_0A92_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a179_1 ( .OUT(na179_1), .IN1(1'b1), .IN2(~na180_1), .IN3(na185_2), .IN4(1'b1), .IN5(na1653_2), .IN6(1'b1), .IN7(1'b0), .IN8(na184_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x37y76     80'h00_0018_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a180_1 ( .OUT(na180_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na40_1), .IN6(~na1025_1), .IN7(1'b0), .IN8(na181_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x46y66     80'h00_0018_00_0000_0CEE_C500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a181_1 ( .OUT(na181_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na431_1), .IN6(1'b0), .IN7(1'b0), .IN8(na164_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x50y58     80'h00_0018_00_0000_0666_F5EC
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a182_1 ( .OUT(na182_1), .IN1(1'b1), .IN2(~na166_1), .IN3(~na868_1), .IN4(~na90_1), .IN5(na908_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x48y70     80'h00_0018_00_0040_0C76_3C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a184_1 ( .OUT(na184_1), .IN1(1'b1), .IN2(~na1813_2), .IN3(~na1593_2), .IN4(1'b0), .IN5(1'b1), .IN6(na893_2), .IN7(1'b1),
                     .IN8(~na39_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x50y73     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a185_4 ( .OUT(na185_2), .IN1(na931_1), .IN2(1'b0), .IN3(na726_2), .IN4(na1594_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x39y71     80'h00_0018_00_0000_0666_09C9
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a186_1 ( .OUT(na186_1), .IN1(na187_1), .IN2(~na191_2), .IN3(1'b0), .IN4(na190_1), .IN5(na189_2), .IN6(~na41_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x37y71     80'h00_0018_00_0040_0C49_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a187_1 ( .OUT(na187_1), .IN1(na40_1), .IN2(1'b0), .IN3(1'b1), .IN4(na1628_2), .IN5(1'b1), .IN6(na1025_1), .IN7(1'b1), .IN8(na181_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x40y72     80'h00_0018_00_0000_0C66_C900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a188_1 ( .OUT(na188_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na189_2), .IN6(~na41_1), .IN7(1'b0), .IN8(na190_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x49y67     80'h00_0060_00_0000_0C0E_FF0D
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a189_4 ( .OUT(na189_2), .IN1(~na431_1), .IN2(na1079_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x34y72     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a190_1 ( .OUT(na190_1), .IN1(1'b1), .IN2(na875_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na616_1), .IN8(~na1026_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x49y72     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a191_4 ( .OUT(na191_2), .IN1(na895_2), .IN2(na727_1), .IN3(1'b0), .IN4(na1594_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x52y74     80'h00_0018_00_0040_0A9B_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a192_1 ( .OUT(na192_1), .IN1(~na1709_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1594_1), .IN5(~na931_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(~na1758_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x48y67     80'h00_0018_00_0040_0C16_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a193_1 ( .OUT(na193_1), .IN1(1'b1), .IN2(na1657_2), .IN3(na195_1), .IN4(1'b0), .IN5(na194_1), .IN6(1'b1), .IN7(1'b1), .IN8(na201_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x45y71     80'h00_0018_00_0040_0C76_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a194_1 ( .OUT(na194_1), .IN1(1'b1), .IN2(~na191_2), .IN3(~na1655_2), .IN4(1'b0), .IN5(~na187_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na188_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x44y71     80'h00_0018_00_0000_0666_9306
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a195_1 ( .OUT(na195_1), .IN1(na199_1), .IN2(na196_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na200_2), .IN7(na198_1),
                     .IN8(~na42_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x35y68     80'h00_0018_00_0040_0C86_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a196_1 ( .OUT(na196_1), .IN1(1'b0), .IN2(na41_1), .IN3(na1629_2), .IN4(1'b1), .IN5(na189_2), .IN6(1'b1), .IN7(1'b1), .IN8(na190_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x34y71     80'h00_0018_00_0000_0C66_9A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a197_1 ( .OUT(na197_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na199_1), .IN6(1'b0), .IN7(na198_1), .IN8(~na42_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x46y63     80'h00_0018_00_0000_0CEE_A500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a198_1 ( .OUT(na198_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na431_1), .IN6(1'b0), .IN7(na1080_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x33y71     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a199_1 ( .OUT(na199_1), .IN1(1'b1), .IN2(na875_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na616_2), .IN8(~na1027_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x49y70     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a200_4 ( .OUT(na200_2), .IN1(1'b0), .IN2(na728_1), .IN3(na1595_1), .IN4(na933_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x52y68     80'h00_0018_00_0040_0A9B_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a201_1 ( .OUT(na201_1), .IN1(1'b1), .IN2(~na727_1), .IN3(1'b1), .IN4(na1594_2), .IN5(~na895_2), .IN6(1'b1), .IN7(1'b0), .IN8(~na1751_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x50y69     80'h00_0018_00_0040_0C16_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a202_1 ( .OUT(na202_1), .IN1(1'b1), .IN2(na204_1), .IN3(na1659_2), .IN4(1'b0), .IN5(na203_1), .IN6(1'b1), .IN7(na210_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x47y67     80'h00_0018_00_0040_0C76_A300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a203_1 ( .OUT(na203_1), .IN1(1'b1), .IN2(~na200_2), .IN3(~na1658_2), .IN4(1'b0), .IN5(1'b1), .IN6(~na196_1), .IN7(na197_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x35y70     80'h00_0018_00_0000_0666_9A3A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a204_1 ( .OUT(na204_1), .IN1(na205_1), .IN2(1'b0), .IN3(1'b0), .IN4(~na209_2), .IN5(na207_2), .IN6(1'b0), .IN7(~na43_1),
                     .IN8(na208_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x35y69     80'h00_0018_00_0040_0C49_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a205_1 ( .OUT(na205_1), .IN1(na1630_2), .IN2(1'b0), .IN3(1'b1), .IN4(na42_1), .IN5(~na199_1), .IN6(1'b1), .IN7(na198_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x36y72     80'h00_0018_00_0000_0C66_9A00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a206_1 ( .OUT(na206_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na207_2), .IN6(1'b0), .IN7(~na43_1), .IN8(na208_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x51y69     80'h00_0060_00_0000_0C0E_FFC5
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a207_4 ( .OUT(na207_2), .IN1(~na431_1), .IN2(1'b0), .IN3(1'b0), .IN4(na1081_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x36y70     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a208_1 ( .OUT(na208_1), .IN1(1'b1), .IN2(~na875_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1028_1), .IN8(~na618_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x52y70     80'h00_0060_00_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a209_4 ( .OUT(na209_2), .IN1(na897_2), .IN2(na729_1), .IN3(na1595_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y69     80'h00_0018_00_0040_0A9B_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a210_1 ( .OUT(na210_1), .IN1(1'b1), .IN2(~na728_1), .IN3(na1595_1), .IN4(1'b1), .IN5(~na1759_2), .IN6(1'b1), .IN7(1'b0),
                     .IN8(~na933_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y64     80'h00_0018_00_0040_0A61_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a211_1 ( .OUT(na211_1), .IN1(na212_1), .IN2(1'b1), .IN3(na219_1), .IN4(1'b1), .IN5(1'b1), .IN6(na213_1), .IN7(na1661_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x39y77     80'h00_0018_00_0040_0CB9_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a212_1 ( .OUT(na212_1), .IN1(~na1660_2), .IN2(1'b1), .IN3(1'b0), .IN4(~na209_2), .IN5(na205_1), .IN6(1'b1), .IN7(1'b1), .IN8(na206_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x39y76     80'h00_0018_00_0000_0666_39CA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a213_1 ( .OUT(na213_1), .IN1(na214_1), .IN2(1'b0), .IN3(1'b0), .IN4(na217_1), .IN5(~na44_1), .IN6(na216_1), .IN7(1'b0), .IN8(~na218_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x39y73     80'h00_0018_00_0040_0A68_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a214_1 ( .OUT(na214_1), .IN1(na207_2), .IN2(1'b1), .IN3(1'b1), .IN4(na208_1), .IN5(1'b0), .IN6(na1631_2), .IN7(na43_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x38y72     80'h00_0018_00_0000_0C66_C900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a215_1 ( .OUT(na215_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na44_1), .IN6(na216_1), .IN7(1'b0), .IN8(na217_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x47y64     80'h00_0018_00_0000_0CEE_A500
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a216_1 ( .OUT(na216_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na431_1), .IN6(1'b0), .IN7(na1082_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x32y72     80'h00_0018_00_0040_0ACC_00F3
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a217_1 ( .OUT(na217_1), .IN1(1'b1), .IN2(~na875_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1029_2), .IN8(~na618_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x44y70     80'h00_0060_00_0000_0C06_FFC6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a218_4 ( .OUT(na218_2), .IN1(na730_1), .IN2(na935_2), .IN3(1'b0), .IN4(na1596_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x52y77     80'h00_0018_00_0040_0A9B_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a219_1 ( .OUT(na219_1), .IN1(1'b1), .IN2(~na729_1), .IN3(na1595_2), .IN4(1'b1), .IN5(~na897_2), .IN6(1'b1), .IN7(1'b0), .IN8(~na1753_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x44y77     80'h00_0018_00_0040_0A92_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a220_1 ( .OUT(na220_1), .IN1(1'b1), .IN2(~na221_1), .IN3(1'b1), .IN4(na228_1), .IN5(na222_1), .IN6(1'b1), .IN7(1'b0), .IN8(na1663_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x47y70     80'h00_0018_00_0040_0CB9_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a221_1 ( .OUT(na221_1), .IN1(~na1662_2), .IN2(1'b1), .IN3(1'b0), .IN4(~na218_2), .IN5(na214_1), .IN6(1'b1), .IN7(1'b1), .IN8(na215_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x39y75     80'h00_0018_00_0000_0666_099A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a222_1 ( .OUT(na222_1), .IN1(na223_1), .IN2(1'b0), .IN3(~na227_2), .IN4(na226_1), .IN5(~na45_1), .IN6(na225_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x33y67     80'h00_0018_00_0040_0C49_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a223_1 ( .OUT(na223_1), .IN1(na44_1), .IN2(1'b0), .IN3(1'b1), .IN4(na1632_2), .IN5(1'b1), .IN6(~na216_1), .IN7(1'b1), .IN8(na217_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x38y74     80'h00_0018_00_0000_0C66_C900
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a224_1 ( .OUT(na224_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na45_1), .IN6(na225_2), .IN7(1'b0), .IN8(na226_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x47y64     80'h00_0060_00_0000_0C0E_FF0B
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a225_4 ( .OUT(na225_2), .IN1(na1083_1), .IN2(~na1674_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x34y74     80'h00_0018_00_0040_0ACC_00FC
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a226_1 ( .OUT(na226_1), .IN1(1'b1), .IN2(na875_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na620_1), .IN8(~na1030_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x42y75     80'h00_0060_00_0000_0C06_FF6C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a227_4 ( .OUT(na227_2), .IN1(1'b0), .IN2(na899_2), .IN3(na731_1), .IN4(na1596_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x44y78     80'h00_0018_00_0040_0C76_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a228_1 ( .OUT(na228_1), .IN1(1'b1), .IN2(~na935_2), .IN3(~na1760_2), .IN4(1'b0), .IN5(na730_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1596_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x46y67     80'h00_0018_00_0040_0A61_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a229_1 ( .OUT(na229_1), .IN1(na230_1), .IN2(1'b1), .IN3(na237_1), .IN4(1'b1), .IN5(1'b1), .IN6(na231_1), .IN7(na1665_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x43y75     80'h00_0018_00_0040_0C76_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a230_1 ( .OUT(na230_1), .IN1(1'b1), .IN2(~na1664_2), .IN3(~na227_2), .IN4(1'b0), .IN5(~na223_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na224_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x41y74     80'h00_0018_00_0000_0666_9C09
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a231_1 ( .OUT(na231_1), .IN1(~na236_2), .IN2(na232_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na234_2), .IN7(~na46_1),
                     .IN8(na235_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x41y78     80'h00_0018_00_0040_0C49_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a232_1 ( .OUT(na232_1), .IN1(na45_1), .IN2(1'b0), .IN3(1'b1), .IN4(na1633_2), .IN5(1'b1), .IN6(~na225_2), .IN7(1'b1), .IN8(na226_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x44y74     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a233_1 ( .OUT(na233_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na234_2), .IN7(~na46_1), .IN8(na235_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x37y72     80'h00_0060_00_0000_0C0E_FF0D
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a234_4 ( .OUT(na234_2), .IN1(~na431_1), .IN2(na1084_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x36y78     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a235_1 ( .OUT(na235_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na875_2), .IN7(1'b1), .IN8(~na1052_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x41y75     80'h00_0060_00_0000_0C06_FF6A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a236_4 ( .OUT(na236_2), .IN1(na937_1), .IN2(1'b0), .IN3(na1597_1), .IN4(na732_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x54y79     80'h00_0018_00_0040_0C76_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a237_1 ( .OUT(na237_1), .IN1(1'b1), .IN2(~na899_2), .IN3(~na1755_2), .IN4(1'b0), .IN5(na1715_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na1596_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x40y75     80'h00_0018_00_0040_0C16_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a238_1 ( .OUT(na238_1), .IN1(1'b1), .IN2(na240_1), .IN3(na1667_2), .IN4(1'b0), .IN5(na239_1), .IN6(1'b1), .IN7(na243_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x41y77     80'h00_0018_00_0040_0CB9_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a239_1 ( .OUT(na239_1), .IN1(~na236_2), .IN2(1'b1), .IN3(1'b0), .IN4(~na1666_2), .IN5(1'b1), .IN6(na232_1), .IN7(1'b1), .IN8(na233_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x41y76     80'h00_0018_00_0000_0666_096C
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a240_1 ( .OUT(na240_1), .IN1(1'b0), .IN2(na1085_1), .IN3(na1597_2), .IN4(na733_1), .IN5(~na47_1), .IN6(na901_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x37y76     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a241_4 ( .OUT(na241_2), .IN1(~na47_1), .IN2(na1085_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x53y81     80'h00_0018_00_0000_0C66_6C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a242_1 ( .OUT(na242_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na901_2), .IN7(na1597_2), .IN8(na733_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x44y79     80'h00_0018_00_0040_0CB9_A300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a243_1 ( .OUT(na243_1), .IN1(~na937_1), .IN2(1'b1), .IN3(1'b0), .IN4(~na1761_2), .IN5(1'b1), .IN6(~na1718_2), .IN7(na1597_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x44y75     80'h00_0018_00_0040_0C29_A300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a244_1 ( .OUT(na244_1), .IN1(na247_1), .IN2(1'b1), .IN3(1'b0), .IN4(na1668_2), .IN5(1'b1), .IN6(~na245_2), .IN7(na250_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ORAND/      x43y76     80'h00_0060_00_0000_0C08_FF37
C_ORAND    #(.CPE_CFG (9'b0_1000_0000)) 
           _a245_4 ( .OUT(na245_2), .IN1(~na242_1), .IN2(~na241_2), .IN3(1'b0), .IN4(~na246_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x38y76     80'h00_0018_00_0040_0A71_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a246_1 ( .OUT(na246_1), .IN1(1'b1), .IN2(na234_2), .IN3(1'b1), .IN4(na235_1), .IN5(~na47_1), .IN6(na1087_1), .IN7(na1803_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x43y77     80'h00_0018_00_0000_0666_9ACA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a247_1 ( .OUT(na247_1), .IN1(na734_2), .IN2(1'b0), .IN3(1'b0), .IN4(na1088_1), .IN5(na734_1), .IN6(1'b0), .IN7(~na48_1),
                     .IN8(na1598_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x33y76     80'h00_0060_00_0000_0C06_FF90
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a248_4 ( .OUT(na248_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na48_1), .IN4(na1088_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x51y81     80'h00_0018_00_0000_0C66_C600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a249_1 ( .OUT(na249_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na734_1), .IN6(na1722_2), .IN7(1'b0), .IN8(na1598_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x56y79     80'h00_0018_00_0040_0A67_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a250_1 ( .OUT(na250_1), .IN1(na1719_2), .IN2(1'b1), .IN3(na1597_2), .IN4(1'b1), .IN5(1'b1), .IN6(~na901_2), .IN7(~na1757_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////D      x47y63     80'h00_FE18_00_0000_0666_60AA
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a251_1 ( .OUT(na251_1), .IN1(na1075_1), .IN2(1'b0), .IN3(na177_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na721_1), .IN8(~na176_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a251_5 ( .OUT(na251_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na251_1) );
// C_XOR///XOR/      x49y66     80'h00_0078_00_0000_0C66_6A63
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a252_1 ( .OUT(na252_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na186_1), .IN6(1'b0), .IN7(na179_1), .IN8(na192_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a252_4 ( .OUT(na252_2), .IN1(1'b0), .IN2(~na284_1), .IN3(na285_2), .IN4(na725_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x49y65     80'h00_0078_00_0000_0C66_A66A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a254_1 ( .OUT(na254_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na203_1), .IN6(na204_1), .IN7(na210_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a254_4 ( .OUT(na254_2), .IN1(na194_1), .IN2(1'b0), .IN3(na195_1), .IN4(na201_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x51y67     80'h00_0078_00_0000_0C66_C6A6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a256_1 ( .OUT(na256_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na222_1), .IN6(na221_1), .IN7(1'b0), .IN8(na228_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a256_4 ( .OUT(na256_2), .IN1(na212_1), .IN2(na213_1), .IN3(na219_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x51y61     80'h00_0078_00_0000_0C66_A6A6
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a258_1 ( .OUT(na258_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na239_1), .IN6(na240_1), .IN7(na243_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a258_4 ( .OUT(na258_2), .IN1(na230_1), .IN2(na231_1), .IN3(na237_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x53y66     80'h00_0060_00_0000_0C06_FFA6
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a259_4 ( .OUT(na259_2), .IN1(na247_1), .IN2(na245_2), .IN3(na250_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x39y79     80'h00_0018_00_0000_0666_999A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a260_1 ( .OUT(na260_1), .IN1(na49_1), .IN2(1'b0), .IN3(na261_1), .IN4(~na265_1), .IN5(na735_1), .IN6(~na1814_2), .IN7(~na940_2),
                     .IN8(na1091_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ORAND////      x44y73     80'h00_0018_00_0000_0C88_37FF
C_ORAND    #(.CPE_CFG (9'b0_0000_0000)) 
           _a261_1 ( .OUT(na261_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na249_1), .IN6(~na248_2), .IN7(1'b0), .IN8(~na262_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x36y76     80'h00_0018_00_0040_0AD4_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a262_1 ( .OUT(na262_1), .IN1(1'b1), .IN2(na234_2), .IN3(1'b1), .IN4(~na235_1), .IN5(na1090_2), .IN6(1'b0), .IN7(~na48_1),
                     .IN8(na1804_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x52y82     80'h00_0018_00_0040_0A9B_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a265_1 ( .OUT(na265_1), .IN1(~na734_1), .IN2(1'b1), .IN3(1'b1), .IN4(na1598_1), .IN5(~na734_2), .IN6(1'b1), .IN7(1'b0), .IN8(~na1723_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y67     80'h00_0018_00_0040_0A92_00A5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a267_1 ( .OUT(na267_1), .IN1(~na1651_2), .IN2(1'b1), .IN3(na721_1), .IN4(1'b1), .IN5(na1075_1), .IN6(1'b1), .IN7(1'b0), .IN8(na1801_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x51y64     80'h00_0018_00_0040_0CD9_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a269_1 ( .OUT(na269_1), .IN1(~na1578_2), .IN2(1'b0), .IN3(1'b1), .IN4(~na1809_2), .IN5(1'b1), .IN6(na889_2), .IN7(1'b1),
                     .IN8(na35_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x47y66     80'h00_0018_00_0040_0CB9_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a272_1 ( .OUT(na272_1), .IN1(~na722_2), .IN2(1'b1), .IN3(1'b0), .IN4(~na1704_2), .IN5(1'b1), .IN6(na269_1), .IN7(1'b1), .IN8(na176_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x37y77     80'h00_0018_00_0040_0CB9_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a274_1 ( .OUT(na274_1), .IN1(~na1810_2), .IN2(1'b1), .IN3(1'b0), .IN4(~na1592_1), .IN5(na36_1), .IN6(1'b1), .IN7(na927_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x52y63     80'h00_0078_00_0000_0C66_369A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a275_1 ( .OUT(na275_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na37_1), .IN6(na891_2), .IN7(1'b0), .IN8(~na1592_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a275_4 ( .OUT(na275_2), .IN1(na38_1), .IN2(1'b0), .IN3(~na1593_1), .IN4(na929_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x53y62     80'h00_0018_00_0040_0CB9_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a277_1 ( .OUT(na277_1), .IN1(~na1705_2), .IN2(1'b1), .IN3(1'b0), .IN4(~na723_1), .IN5(na274_1), .IN6(1'b1), .IN7(na275_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x35y72     80'h00_0018_00_0040_0CB9_CA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a279_1 ( .OUT(na279_1), .IN1(~na1811_2), .IN2(1'b1), .IN3(1'b0), .IN4(~na1592_2), .IN5(na37_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1748_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x53y61     80'h00_0018_00_0040_0CB9_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a282_1 ( .OUT(na282_1), .IN1(~na724_1), .IN2(1'b1), .IN3(1'b0), .IN4(~na1706_2), .IN5(1'b1), .IN6(na279_1), .IN7(na275_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x37y78     80'h00_0018_00_0040_0C76_C500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a284_1 ( .OUT(na284_1), .IN1(1'b1), .IN2(~na1812_2), .IN3(~na1593_1), .IN4(1'b0), .IN5(~na38_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na929_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x52y71     80'h00_0060_00_0000_0C06_FF9C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a285_4 ( .OUT(na285_2), .IN1(1'b0), .IN2(na893_2), .IN3(~na1593_2), .IN4(na39_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x54y63     80'h00_0018_00_0040_0CB9_AC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a288_1 ( .OUT(na288_1), .IN1(~na1707_2), .IN2(1'b1), .IN3(1'b0), .IN4(~na725_1), .IN5(1'b1), .IN6(na284_1), .IN7(na285_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x49y61     80'h00_0078_00_0000_0C66_9966
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a290_1 ( .OUT(na290_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na274_1), .IN6(na272_1), .IN7(na275_1), .IN8(~na723_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a290_4 ( .OUT(na290_2), .IN1(~na722_2), .IN2(~na269_1), .IN3(na267_1), .IN4(na176_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x52y64     80'h00_0078_00_0000_0C66_9999
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a292_1 ( .OUT(na292_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na282_1), .IN6(~na284_1), .IN7(na285_2), .IN8(~na725_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a292_4 ( .OUT(na292_2), .IN1(~na724_1), .IN2(na277_1), .IN3(na275_2), .IN4(~na1670_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x48y63     80'h00_0018_00_0000_0666_6660
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a293_1 ( .OUT(na293_1), .IN1(1'b0), .IN2(1'b0), .IN3(na288_1), .IN4(na184_1), .IN5(~na40_1), .IN6(~na1025_1), .IN7(~na185_2),
                     .IN8(~na181_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x55y76     80'h00_0018_00_0040_0C16_AA00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a295_1 ( .OUT(na295_1), .IN1(1'b1), .IN2(na901_1), .IN3(na1756_2), .IN4(1'b0), .IN5(na897_1), .IN6(1'b1), .IN7(na108_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x57y79     80'h00_0018_00_0000_0C88_65FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a296_1 ( .OUT(na296_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1100_1), .IN6(1'b0), .IN7(na1754_2), .IN8(~na963_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x58y79     80'h00_0018_00_0040_0C42_3300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a297_1 ( .OUT(na297_1), .IN1(1'b0), .IN2(na899_1), .IN3(1'b1), .IN4(1'b0), .IN5(1'b1), .IN6(~na1772_2), .IN7(1'b1), .IN8(~na963_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x53y79     80'h00_0018_00_0040_0C18_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a298_1 ( .OUT(na298_1), .IN1(1'b1), .IN2(1'b0), .IN3(1'b0), .IN4(na960_1), .IN5(1'b1), .IN6(~na901_1), .IN7(1'b1), .IN8(na963_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x53y82     80'h00_0018_00_0040_0C42_3500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a299_1 ( .OUT(na299_1), .IN1(1'b0), .IN2(na901_1), .IN3(1'b1), .IN4(1'b0), .IN5(~na1773_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na963_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x58y72     80'h00_0018_00_0040_0C49_5C00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a300_1 ( .OUT(na300_1), .IN1(na303_1), .IN2(1'b0), .IN3(1'b1), .IN4(na1672_2), .IN5(1'b1), .IN6(na893_1), .IN7(~na301_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x58y73     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a301_1 ( .OUT(na301_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na302_2), .IN8(na963_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x60y73     80'h00_0060_00_0000_0C08_FF11
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a302_4 ( .OUT(na302_2), .IN1(~na1747_2), .IN2(~na891_1), .IN3(~na965_1), .IN4(~na957_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x55y69     80'h00_0018_00_0000_0C66_9C00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a303_1 ( .OUT(na303_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1778_2), .IN7(~na119_2), .IN8(na957_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x54y69     80'h00_0060_00_0000_0C08_FFC6
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a304_4 ( .OUT(na304_2), .IN1(na1647_2), .IN2(~na889_1), .IN3(1'b0), .IN4(~na121_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x56y72     80'h00_0018_00_0000_0CEE_CE00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a305_1 ( .OUT(na305_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1647_2), .IN6(na889_1), .IN7(1'b0), .IN8(na1102_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x57y72     80'h00_0078_00_0000_0CEE_A53C
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a307_1 ( .OUT(na307_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1061_1), .IN6(1'b0), .IN7(na127_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a307_4 ( .OUT(na307_2), .IN1(1'b0), .IN2(na125_2), .IN3(1'b0), .IN4(~na1060_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x58y69     80'h00_0078_00_0000_0CEE_A3C5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a309_1 ( .OUT(na309_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(~na1063_1), .IN7(na131_1), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a309_4 ( .OUT(na309_2), .IN1(~na1062_1), .IN2(1'b0), .IN3(1'b0), .IN4(na129_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x58y76     80'h00_0078_00_0000_0CEE_0DA5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a311_1 ( .OUT(na311_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1065_1), .IN6(na135_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a311_4 ( .OUT(na311_2), .IN1(~na1064_1), .IN2(1'b0), .IN3(na133_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x60y77     80'h00_0060_00_0000_0C0E_FFC5
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a312_4 ( .OUT(na312_2), .IN1(~na1066_1), .IN2(1'b0), .IN3(1'b0), .IN4(na137_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x56y78     80'h00_0018_00_0000_0666_3FBC
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a314_1 ( .OUT(na314_1), .IN1(1'b1), .IN2(~na899_1), .IN3(~na958_1), .IN4(na1774_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na963_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x56y81     80'h00_0018_00_0000_0C88_4FFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a318_1 ( .OUT(na318_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(~na962_1), .IN8(na963_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x60y75     80'h00_0018_00_0000_0666_F3B5
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a319_1 ( .OUT(na319_1), .IN1(na303_1), .IN2(1'b1), .IN3(~na302_2), .IN4(na963_1), .IN5(1'b1), .IN6(na893_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x56y70     80'h00_0018_00_0040_0C29_A300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a321_1 ( .OUT(na321_1), .IN1(na1720_2), .IN2(1'b1), .IN3(1'b0), .IN4(na733_2), .IN5(1'b1), .IN6(~na729_2), .IN7(na108_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x60y79     80'h00_0060_00_0000_0C08_FF36
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a322_4 ( .OUT(na322_2), .IN1(na1716_2), .IN2(~na979_1), .IN3(1'b0), .IN4(na1116_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x59y74     80'h00_0018_00_0040_0C24_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a323_1 ( .OUT(na323_1), .IN1(1'b0), .IN2(1'b1), .IN3(na731_2), .IN4(1'b0), .IN5(1'b1), .IN6(na976_1), .IN7(1'b1), .IN8(na1791_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x62y77     80'h00_0018_00_0040_0C42_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a324_1 ( .OUT(na324_1), .IN1(1'b0), .IN2(na976_1), .IN3(1'b1), .IN4(1'b0), .IN5(1'b1), .IN6(na979_1), .IN7(1'b1), .IN8(na733_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x54y81     80'h00_0018_00_0040_0C18_A500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a325_1 ( .OUT(na325_1), .IN1(1'b1), .IN2(1'b0), .IN3(1'b0), .IN4(na733_2), .IN5(~na978_1), .IN6(1'b1), .IN7(na1790_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x48y65     80'h00_0018_00_0040_0C16_CC00
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a326_1 ( .OUT(na326_1), .IN1(1'b1), .IN2(na329_1), .IN3(na1673_2), .IN4(1'b0), .IN5(1'b1), .IN6(na327_2), .IN7(1'b1), .IN8(na725_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x55y68     80'h00_0060_00_0000_0C08_FFF4
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a327_4 ( .OUT(na327_2), .IN1(~na328_1), .IN2(na979_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x53y63     80'h00_0018_00_0000_0C88_11FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a328_1 ( .OUT(na328_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na981_1), .IN6(~na973_1), .IN7(~na721_2), .IN8(~na723_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x55y68     80'h00_0018_00_0000_0C66_5600
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a329_1 ( .OUT(na329_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1793_2), .IN6(na973_1), .IN7(~na119_2), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x54y67     80'h00_0060_00_0000_0C08_FF6C
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a330_4 ( .OUT(na330_2), .IN1(1'b0), .IN2(~na139_1), .IN3(~na721_2), .IN4(na116_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR////      x53y66     80'h00_0018_00_0000_0CEE_EC00
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a331_1 ( .OUT(na331_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1118_2), .IN7(na721_2), .IN8(na116_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x58y65     80'h00_0078_00_0000_0CEE_0DD0
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a333_1 ( .OUT(na333_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na1068_1), .IN6(na145_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a333_4 ( .OUT(na333_2), .IN1(1'b0), .IN2(1'b0), .IN3(~na1067_1), .IN4(na143_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x59y69     80'h00_0078_00_0000_0CEE_0BA5
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a335_1 ( .OUT(na335_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na149_2), .IN6(~na1070_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a335_4 ( .OUT(na335_2), .IN1(~na1069_1), .IN2(1'b0), .IN3(na147_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_OR///OR/      x58y75     80'h00_0078_00_0000_0CEE_B00D
C_OR       #(.CPE_CFG (9'b0_0000_0000)) 
           _a337_1 ( .OUT(na337_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na153_2), .IN8(~na1072_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a337_4 ( .OUT(na337_2), .IN1(~na1071_1), .IN2(na151_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///OR/      x58y71     80'h00_0060_00_0000_0C0E_FFA5
C_OR       #(.CPE_CFG (9'b0_1000_0000)) 
           _a338_4 ( .OUT(na338_2), .IN1(~na1073_1), .IN2(1'b0), .IN3(na155_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x53y78     80'h00_0018_00_0000_0666_F3AB
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a340_1 ( .OUT(na340_1), .IN1(~na974_1), .IN2(na1788_2), .IN3(~na731_2), .IN4(1'b1), .IN5(1'b1), .IN6(na979_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x55y80     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a344_1 ( .OUT(na344_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na978_1), .IN6(na979_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ANDXOR////      x47y65     80'h00_0018_00_0000_0666_3F5B
C_ANDXOR   #(.CPE_CFG (9'b0_0000_0000)) 
           _a345_1 ( .OUT(na345_1), .IN1(~na328_1), .IN2(na979_1), .IN3(na1673_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na725_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x45y66     80'h00_0078_00_0020_0C66_0305
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a411_1 ( .OUT(na411_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na942_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na424_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a411_4 ( .OUT(na411_2), .COUTY1(na411_4), .IN1(~na944_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na942_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na424_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x45y67     80'h00_0018_00_0010_0666_0005
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a413_1 ( .OUT(na413_1), .COUTY1(na413_4), .IN1(~na944_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na411_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////Carry      x45y68     80'h00_0058_00_0010_0666_0003
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a414_1 ( .OUT(na414_1), .COUTY1(na414_4), .IN1(1'b1), .IN2(~na946_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na413_4), .PINX(1'b0), .PINY1(1'b0) );
C_Carry    #(.CPE_CFG (9'bX_0000_0010)) 
           _a414_5 ( .OUT(na414_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(na414_4), .D_IN(na414_1) );
// C_ADDF////      x45y69     80'h00_0018_00_0010_0666_0003
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a415_1 ( .OUT(na415_1), .COUTY1(na415_4), .IN1(1'b1), .IN2(~na946_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na414_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x45y61     80'h00_0078_00_0020_0C66_3503
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a416_1 ( .OUT(na416_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na251_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na173_1),
                     .CINX(1'b0), .CINY1(na425_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a416_4 ( .OUT(na416_2), .COUTY1(na416_4), .IN1(1'b1), .IN2(~na949_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na251_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(~na173_1), .CINX(1'b0), .CINY1(na425_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x45y62     80'h00_0078_00_0020_0C66_0305
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a418_1 ( .OUT(na418_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na949_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na416_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a418_4 ( .OUT(na418_2), .COUTY1(na418_4), .IN1(~na951_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na949_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na416_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x45y63     80'h00_0078_00_0020_0C66_0503
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a420_1 ( .OUT(na420_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na951_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na418_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a420_4 ( .OUT(na420_2), .COUTY1(na420_4), .IN1(1'b1), .IN2(~na953_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na951_2), .IN6(1'b1),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na418_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x45y64     80'h00_0078_00_0020_0C66_0305
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a422_1 ( .OUT(na422_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na953_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na420_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a422_4 ( .OUT(na422_2), .COUTY1(na422_4), .IN1(~na955_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na953_2),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na420_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x45y65     80'h00_0078_00_0020_0C66_0503
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a424_1 ( .OUT(na424_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na955_2), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na422_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a424_4 ( .OUT(na424_2), .COUTY1(na424_4), .IN1(1'b1), .IN2(~na942_1), .IN3(1'b0), .IN4(1'b0), .IN5(~na955_2), .IN6(1'b1),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na422_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x45y60     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a425_2 ( .OUT(na425_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a425_6 ( .COUTY1(na425_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na425_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x22y67     80'h00_FA60_00_0020_0C66_ACCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a426_1 ( .OUT(na426_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na1738_2), .IN7(na426_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na428_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a426_2 ( .OUT(na426_1), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na426_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a426_4 ( .OUT(na426_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na862_1), .IN5(1'b1), .IN6(na1738_2), .IN7(na426_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na428_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x22y66     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a428_2 ( .OUT(na428_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a428_6 ( .COUTY1(na428_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na428_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x45y58     80'h00_FA60_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a429_1 ( .OUT(na429_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na429_1), .IN7(na904_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na433_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0000)) 
           _a429_2 ( .OUT(na429_1), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na429_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a429_4 ( .OUT(na429_2), .COUTY1(na429_4), .IN1(1'b0), .IN2(1'b0), .IN3(na906_2), .IN4(1'b1), .IN5(1'b1), .IN6(na429_1), .IN7(na904_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na433_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x45y59     80'h00_FA60_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a431_1 ( .OUT(na431_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na431_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na429_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a431_2 ( .OUT(na431_1), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na431_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a431_4 ( .OUT(na431_2), .IN1(na908_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na431_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na429_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x45y57     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a433_2 ( .OUT(na433_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a433_6 ( .COUTY1(na433_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na433_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x48y59     80'h00_0078_00_0020_0C66_AC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a434_1 ( .OUT(na434_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na745_2), .IN7(na744_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na437_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a434_4 ( .OUT(na434_2), .COUTY1(na434_4), .IN1(1'b1), .IN2(na745_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na745_2), .IN7(na744_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na437_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////D      x48y60     80'h00_FE18_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a436_1 ( .OUT(na436_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na436_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na434_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a436_5 ( .OUT(na436_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na436_1) );
// C_/C_0_1///      x48y58     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a437_2 ( .OUT(na437_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a437_6 ( .COUTY1(na437_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na437_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x31y70     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a439_1 ( .OUT(na439_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na45_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na452_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a439_4 ( .OUT(na439_2), .COUTY1(na439_4), .IN1(1'b0), .IN2(1'b0), .IN3(na46_1), .IN4(1'b1), .IN5(na45_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na452_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x31y71     80'h00_0078_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a441_1 ( .OUT(na441_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na47_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na439_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a441_4 ( .OUT(na441_2), .COUTY1(na441_4), .IN1(1'b0), .IN2(1'b0), .IN3(na48_1), .IN4(1'b1), .IN5(na47_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na439_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x31y72     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a443_1 ( .OUT(na443_1), .IN1(na49_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na441_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x31y65     80'h00_0078_00_0020_0C66_CC0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a444_1 ( .OUT(na444_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na844_2), .IN7(1'b1), .IN8(na35_1),
                     .CINX(1'b0), .CINY1(na453_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a444_4 ( .OUT(na444_2), .COUTY1(na444_4), .IN1(na36_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na844_2), .IN7(1'b1),
                     .IN8(na35_1), .CINX(1'b0), .CINY1(na453_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x31y66     80'h00_0078_00_0020_0C66_0A0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a446_1 ( .OUT(na446_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na37_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na444_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a446_4 ( .OUT(na446_2), .COUTY1(na446_4), .IN1(na38_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na37_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na444_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x31y67     80'h00_0078_00_0020_0C66_C00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a448_1 ( .OUT(na448_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(na39_1),
                     .CINX(1'b0), .CINY1(na446_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a448_4 ( .OUT(na448_2), .COUTY1(na448_4), .IN1(na40_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1),
                     .IN8(na39_1), .CINX(1'b0), .CINY1(na446_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x31y68     80'h00_0078_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a450_1 ( .OUT(na450_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na41_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na448_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a450_4 ( .OUT(na450_2), .COUTY1(na450_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na42_1), .IN5(1'b1), .IN6(na41_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na448_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x31y69     80'h00_0078_00_0020_0C66_A00A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a452_1 ( .OUT(na452_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na43_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na450_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a452_4 ( .OUT(na452_2), .COUTY1(na452_4), .IN1(na44_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na43_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na450_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x31y64     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a453_2 ( .OUT(na453_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a453_6 ( .COUTY1(na453_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na453_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x30y70     80'h00_0078_00_0020_0C66_FAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a455_1 ( .OUT(na455_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na45_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na468_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a455_4 ( .OUT(na455_2), .COUTY1(na455_4), .IN1(1'b1), .IN2(1'b1), .IN3(na46_1), .IN4(1'b1), .IN5(na45_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na468_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x30y71     80'h00_0078_00_0020_0C66_FAAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a457_1 ( .OUT(na457_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na47_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na455_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a457_4 ( .OUT(na457_2), .COUTY1(na457_4), .IN1(1'b1), .IN2(1'b1), .IN3(na48_1), .IN4(1'b1), .IN5(na47_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na455_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x30y72     80'h00_0018_00_0010_0666_00FA
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a459_1 ( .OUT(na459_1), .IN1(na49_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na457_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x30y65     80'h00_0078_00_0020_0C66_CCFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a460_1 ( .OUT(na460_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na844_2), .IN7(1'b1), .IN8(na35_1),
                     .CINX(1'b0), .CINY1(na469_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a460_4 ( .OUT(na460_2), .COUTY1(na460_4), .IN1(na36_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na844_2), .IN7(1'b1),
                     .IN8(na35_1), .CINX(1'b0), .CINY1(na469_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x30y66     80'h00_0078_00_0020_0C66_FAFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a462_1 ( .OUT(na462_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na37_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na460_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a462_4 ( .OUT(na462_2), .COUTY1(na462_4), .IN1(na38_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na37_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na460_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x30y67     80'h00_0078_00_0020_0C66_CFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a464_1 ( .OUT(na464_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na39_1),
                     .CINX(1'b0), .CINY1(na462_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a464_4 ( .OUT(na464_2), .COUTY1(na464_4), .IN1(na40_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na39_1), .CINX(1'b0), .CINY1(na462_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x30y68     80'h00_0078_00_0020_0C66_FCCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a466_1 ( .OUT(na466_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na41_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na464_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a466_4 ( .OUT(na466_2), .COUTY1(na466_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na42_1), .IN5(1'b1), .IN6(na41_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na464_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x30y69     80'h00_0078_00_0020_0C66_AFFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a468_1 ( .OUT(na468_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(na43_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na466_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a468_4 ( .OUT(na468_2), .COUTY1(na468_4), .IN1(na44_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na43_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na466_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x30y64     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a469_2 ( .OUT(na469_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a469_6 ( .COUTY1(na469_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na469_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x46y53     80'h00_FE60_00_0020_0C66_0CFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a471_1 ( .OUT(na471_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na495_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a471_2 ( .OUT(na471_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na471_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a471_4 ( .OUT(na471_2), .COUTY1(na471_4), .IN1(1'b1), .IN2(na946_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na946_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na495_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y54     80'h00_FE60_00_0020_0C66_FCFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a473_1 ( .OUT(na473_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na471_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a473_2 ( .OUT(na473_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na473_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a473_4 ( .OUT(na473_2), .COUTY1(na473_4), .IN1(1'b1), .IN2(na946_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na946_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na471_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y55     80'h00_FE60_00_0020_0C66_0CFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a475_1 ( .OUT(na475_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na473_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a475_2 ( .OUT(na475_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na475_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a475_4 ( .OUT(na475_2), .COUTY1(na475_4), .IN1(1'b1), .IN2(na946_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na946_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na473_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y56     80'h00_FE60_00_0020_0C66_FC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a477_1 ( .OUT(na477_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na475_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a477_2 ( .OUT(na477_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na477_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a477_4 ( .OUT(na477_2), .COUTY1(na477_4), .IN1(1'b1), .IN2(na946_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na475_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y57     80'h00_FE60_00_0020_0C66_0CFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a479_1 ( .OUT(na479_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na477_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a479_2 ( .OUT(na479_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na479_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a479_4 ( .OUT(na479_2), .COUTY1(na479_4), .IN1(1'b1), .IN2(na946_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na946_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na477_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y48     80'h00_FE60_00_0020_0C66_AA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a480_1 ( .OUT(na480_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na951_1), .IN6(1'b1), .IN7(na1766_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na496_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a480_2 ( .OUT(na480_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na480_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a480_4 ( .OUT(na480_2), .COUTY1(na480_4), .IN1(1'b1), .IN2(na953_1), .IN3(1'b0), .IN4(1'b0), .IN5(na951_1), .IN6(1'b1), .IN7(na1766_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na496_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y58     80'h00_FE60_00_0020_0C66_FC0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a482_1 ( .OUT(na482_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na479_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a482_2 ( .OUT(na482_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na482_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a482_4 ( .OUT(na482_2), .COUTY1(na482_4), .IN1(1'b1), .IN2(na946_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na479_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y59     80'h00_FE60_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a484_1 ( .OUT(na484_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na482_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a484_2 ( .OUT(na484_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na484_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a484_4 ( .OUT(na484_2), .COUTY1(na484_4), .IN1(1'b1), .IN2(na946_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na482_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y60     80'h00_FE60_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a486_1 ( .OUT(na486_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na484_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a486_2 ( .OUT(na486_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na486_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a486_4 ( .OUT(na486_2), .IN1(1'b1), .IN2(na946_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na946_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na484_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y49     80'h00_FE60_00_0020_0C66_0C0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a489_1 ( .OUT(na489_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na953_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na480_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a489_2 ( .OUT(na489_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na489_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a489_4 ( .OUT(na489_2), .COUTY1(na489_4), .IN1(na955_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na953_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na480_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y50     80'h00_FE60_00_0020_0C66_FAFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a491_1 ( .OUT(na491_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na955_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na489_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a491_2 ( .OUT(na491_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na491_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a491_4 ( .OUT(na491_2), .COUTY1(na491_4), .IN1(1'b1), .IN2(na942_1), .IN3(1'b1), .IN4(1'b1), .IN5(na955_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na489_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y51     80'h00_FE60_00_0020_0C66_0CFA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a493_1 ( .OUT(na493_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na942_2), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na491_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a493_2 ( .OUT(na493_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na493_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a493_4 ( .OUT(na493_2), .COUTY1(na493_4), .IN1(na944_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na942_2), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na491_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x46y52     80'h00_FE60_00_0020_0C66_FA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a495_1 ( .OUT(na495_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na944_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na493_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a495_2 ( .OUT(na495_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na495_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a495_4 ( .OUT(na495_2), .COUTY1(na495_4), .IN1(1'b1), .IN2(na946_1), .IN3(1'b0), .IN4(1'b0), .IN5(na944_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na493_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x46y47     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a496_2 ( .OUT(na496_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a496_6 ( .COUTY1(na496_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na496_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x57y65     80'h00_FE60_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a498_1 ( .OUT(na498_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na498_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na511_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a498_2 ( .OUT(na498_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na498_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a498_4 ( .OUT(na498_2), .COUTY1(na498_4), .IN1(1'b0), .IN2(1'b0), .IN3(na706_1), .IN4(1'b1), .IN5(na498_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na511_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x57y66     80'h00_FE60_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a500_1 ( .OUT(na500_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na500_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na498_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a500_2 ( .OUT(na500_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na500_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a500_4 ( .OUT(na500_2), .COUTY1(na500_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na708_2), .IN5(1'b1), .IN6(na500_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na498_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF/D///      x57y67     80'h00_FE00_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a502_1 ( .OUT(na502_1_i), .IN1(na502_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na500_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a502_2 ( .OUT(na502_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na502_1_i) );
// C_ADDF2/D//ADDF2/      x57y60     80'h00_FE60_00_0020_0C66_ACA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a503_1 ( .OUT(na503_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na503_1), .IN7(na696_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na540_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a503_2 ( .OUT(na503_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na503_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a503_4 ( .OUT(na503_2), .COUTY1(na503_4), .IN1(1'b0), .IN2(1'b0), .IN3(na696_1), .IN4(1'b1), .IN5(1'b1), .IN6(na503_1), .IN7(na696_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na540_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x57y61     80'h00_FE60_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a505_1 ( .OUT(na505_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na505_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na503_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a505_2 ( .OUT(na505_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na505_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a505_4 ( .OUT(na505_2), .COUTY1(na505_4), .IN1(1'b0), .IN2(1'b0), .IN3(na698_1), .IN4(1'b1), .IN5(na505_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na503_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x57y62     80'h00_FE60_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a507_1 ( .OUT(na507_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na507_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na505_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a507_2 ( .OUT(na507_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na507_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a507_4 ( .OUT(na507_2), .COUTY1(na507_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na700_2), .IN5(1'b1), .IN6(na507_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na505_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x57y63     80'h00_FE60_00_0020_0C66_0AC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a509_1 ( .OUT(na509_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na509_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na507_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a509_2 ( .OUT(na509_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na509_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a509_4 ( .OUT(na509_2), .COUTY1(na509_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na702_1), .IN5(na509_1), .IN6(1'b1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na507_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x57y64     80'h00_FE60_00_0020_0C66_0CA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a511_1 ( .OUT(na511_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na511_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na509_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a511_2 ( .OUT(na511_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na511_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a511_4 ( .OUT(na511_2), .COUTY1(na511_4), .IN1(1'b0), .IN2(1'b0), .IN3(na704_2), .IN4(1'b1), .IN5(1'b1), .IN6(na511_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na509_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y49     80'h00_FE60_00_0020_0C66_AACC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a512_1 ( .OUT(na512_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1724_2), .IN6(1'b1), .IN7(na512_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na546_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a512_2 ( .OUT(na512_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na512_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a512_4 ( .OUT(na512_2), .COUTY1(na512_4), .IN1(1'b1), .IN2(na776_1), .IN3(1'b1), .IN4(na748_1), .IN5(na1724_2), .IN6(1'b1),
                     .IN7(na512_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na546_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y54     80'h00_FE60_00_0020_0C66_CAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a513_1 ( .OUT(na513_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1729_2), .IN6(1'b1), .IN7(1'b1), .IN8(na513_1),
                     .CINX(1'b0), .CINY1(na538_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a513_2 ( .OUT(na513_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na513_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a513_4 ( .OUT(na513_2), .COUTY1(na513_4), .IN1(na786_1), .IN2(1'b1), .IN3(na758_2), .IN4(1'b1), .IN5(na1729_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na513_1), .CINX(1'b0), .CINY1(na538_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y55     80'h00_FE60_00_0020_0C66_AAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a515_1 ( .OUT(na515_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1730_2), .IN6(1'b1), .IN7(na515_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na513_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a515_2 ( .OUT(na515_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na515_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a515_4 ( .OUT(na515_2), .COUTY1(na515_4), .IN1(1'b1), .IN2(na788_1), .IN3(na760_2), .IN4(1'b1), .IN5(na1730_2), .IN6(1'b1),
                     .IN7(na515_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na513_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y56     80'h00_FE60_00_0020_0C66_CAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a517_1 ( .OUT(na517_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1731_2), .IN6(1'b1), .IN7(1'b1), .IN8(na517_1),
                     .CINX(1'b0), .CINY1(na515_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a517_2 ( .OUT(na517_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na517_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a517_4 ( .OUT(na517_2), .COUTY1(na517_4), .IN1(1'b1), .IN2(na790_1), .IN3(na762_1), .IN4(1'b1), .IN5(na1731_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na517_1), .CINX(1'b0), .CINY1(na515_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y57     80'h00_FE60_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a519_1 ( .OUT(na519_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1732_2), .IN6(1'b1), .IN7(na519_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na517_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a519_2 ( .OUT(na519_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na519_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a519_4 ( .OUT(na519_2), .COUTY1(na519_4), .IN1(na792_1), .IN2(1'b1), .IN3(na764_2), .IN4(1'b1), .IN5(na1732_2), .IN6(1'b1),
                     .IN7(na519_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na517_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y58     80'h00_FE60_00_0020_0C66_CACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a521_1 ( .OUT(na521_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1733_2), .IN6(1'b1), .IN7(1'b1), .IN8(na521_1),
                     .CINX(1'b0), .CINY1(na519_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a521_2 ( .OUT(na521_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na521_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a521_4 ( .OUT(na521_2), .COUTY1(na521_4), .IN1(na766_1), .IN2(1'b1), .IN3(1'b1), .IN4(na794_1), .IN5(na1733_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na521_1), .CINX(1'b0), .CINY1(na519_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y59     80'h00_FE60_00_0020_0C66_AAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a524_1 ( .OUT(na524_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1734_2), .IN6(1'b1), .IN7(na524_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na521_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a524_2 ( .OUT(na524_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na524_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a524_4 ( .OUT(na524_2), .COUTY1(na524_4), .IN1(1'b1), .IN2(na768_1), .IN3(na796_1), .IN4(1'b1), .IN5(na1734_2), .IN6(1'b1),
                     .IN7(na524_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na521_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y60     80'h00_FE60_00_0020_0C66_CAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a526_1 ( .OUT(na526_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1735_2), .IN6(1'b1), .IN7(1'b1), .IN8(na526_1),
                     .CINX(1'b0), .CINY1(na524_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a526_2 ( .OUT(na526_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na526_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a526_4 ( .OUT(na526_2), .COUTY1(na526_4), .IN1(1'b1), .IN2(na798_1), .IN3(na770_1), .IN4(1'b1), .IN5(na1735_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na526_1), .CINX(1'b0), .CINY1(na524_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y61     80'h00_FE60_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a528_1 ( .OUT(na528_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1736_2), .IN6(1'b1), .IN7(na528_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na526_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a528_2 ( .OUT(na528_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na528_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a528_4 ( .OUT(na528_2), .COUTY1(na528_4), .IN1(na800_1), .IN2(1'b1), .IN3(1'b1), .IN4(na772_2), .IN5(na1736_2), .IN6(1'b1),
                     .IN7(na528_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na526_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y62     80'h00_FE60_00_0020_0C66_CAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a530_1 ( .OUT(na530_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1737_2), .IN6(1'b1), .IN7(1'b1), .IN8(na530_1),
                     .CINX(1'b0), .CINY1(na528_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a530_2 ( .OUT(na530_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na530_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a530_4 ( .OUT(na530_2), .IN1(na774_1), .IN2(1'b1), .IN3(na802_1), .IN4(1'b1), .IN5(na1737_2), .IN6(1'b1), .IN7(1'b1), .IN8(na530_1),
                     .CINX(1'b0), .CINY1(na528_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y50     80'h00_FE60_00_0020_0C66_CAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a532_1 ( .OUT(na532_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1725_2), .IN6(1'b1), .IN7(1'b1), .IN8(na532_1),
                     .CINX(1'b0), .CINY1(na512_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a532_2 ( .OUT(na532_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na532_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a532_4 ( .OUT(na532_2), .COUTY1(na532_4), .IN1(1'b1), .IN2(na778_1), .IN3(na750_2), .IN4(1'b1), .IN5(na1725_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na532_1), .CINX(1'b0), .CINY1(na512_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y51     80'h00_FE60_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a534_1 ( .OUT(na534_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1726_2), .IN6(1'b1), .IN7(na534_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na532_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a534_2 ( .OUT(na534_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na534_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a534_4 ( .OUT(na534_2), .COUTY1(na534_4), .IN1(na780_1), .IN2(1'b1), .IN3(na752_1), .IN4(1'b1), .IN5(na1726_2), .IN6(1'b1),
                     .IN7(na534_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na532_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y52     80'h00_FE60_00_0020_0C66_CAAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a536_1 ( .OUT(na536_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1727_2), .IN6(1'b1), .IN7(1'b1), .IN8(na536_1),
                     .CINX(1'b0), .CINY1(na534_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a536_2 ( .OUT(na536_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na536_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a536_4 ( .OUT(na536_2), .COUTY1(na536_4), .IN1(1'b1), .IN2(na782_1), .IN3(na754_1), .IN4(1'b1), .IN5(na1727_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na536_1), .CINX(1'b0), .CINY1(na534_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x52y53     80'h00_FE60_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a538_1 ( .OUT(na538_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1728_2), .IN6(1'b1), .IN7(na538_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na536_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a538_2 ( .OUT(na538_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na538_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a538_4 ( .OUT(na538_2), .COUTY1(na538_4), .IN1(na784_1), .IN2(1'b1), .IN3(na756_2), .IN4(1'b1), .IN5(na1728_2), .IN6(1'b1),
                     .IN7(na538_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na536_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x57y59     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a540_2 ( .OUT(na540_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a540_6 ( .COUTY1(na540_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na540_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x24y77     80'h00_0078_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a541_1 ( .OUT(na541_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na98_2), .IN7(1'b1), .IN8(na99_2),
                     .CINX(1'b0), .CINY1(na552_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a541_4 ( .OUT(na541_2), .COUTY1(na541_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na99_1), .IN5(1'b1), .IN6(na98_2), .IN7(1'b1),
                     .IN8(na99_2), .CINX(1'b0), .CINY1(na552_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x24y78     80'h00_0078_00_0020_0C66_0C0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a543_1 ( .OUT(na543_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na98_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na541_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a543_4 ( .OUT(na543_2), .COUTY1(na543_4), .IN1(na97_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na98_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na541_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x24y79     80'h00_0018_00_0010_0666_00C0
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a545_1 ( .OUT(na545_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na94_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na543_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x52y48     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a546_2 ( .OUT(na546_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a546_6 ( .COUTY1(na546_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na546_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x24y54     80'h00_0078_00_0020_0C66_ACCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a547_1 ( .OUT(na547_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na109_1), .IN7(na110_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na575_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a547_4 ( .OUT(na547_2), .COUTY1(na547_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na107_1), .IN5(1'b1), .IN6(na109_1), .IN7(na110_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na575_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x24y55     80'h00_0078_00_0020_0C66_FAFC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a549_1 ( .OUT(na549_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na106_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na547_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a549_4 ( .OUT(na549_2), .COUTY1(na549_4), .IN1(1'b1), .IN2(na109_2), .IN3(1'b1), .IN4(1'b1), .IN5(na106_2), .IN6(1'b1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na547_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x24y56     80'h00_0018_00_0010_0666_00AF
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a551_1 ( .OUT(na551_1), .IN1(1'b1), .IN2(1'b1), .IN3(na110_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na549_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x24y76     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a552_2 ( .OUT(na552_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a552_6 ( .COUTY1(na552_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na552_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x51y54     80'h00_0078_00_0020_0C66_CA30
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a553_1 ( .OUT(na553_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na165_1), .IN6(1'b1), .IN7(1'b1), .IN8(na164_1),
                     .CINX(1'b0), .CINY1(na581_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a553_4 ( .OUT(na553_2), .COUTY1(na553_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1016_1), .IN5(na165_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na164_1), .CINX(1'b0), .CINY1(na581_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y55     80'h00_0078_00_0020_0C66_0350
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a555_1 ( .OUT(na555_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na1019_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na553_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a555_4 ( .OUT(na555_2), .COUTY1(na555_4), .IN1(1'b0), .IN2(1'b0), .IN3(~na1022_1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1019_1),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na553_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y56     80'h00_0078_00_0020_0C66_30C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a557_1 ( .OUT(na557_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na1024_1),
                     .CINX(1'b0), .CINY1(na555_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a557_4 ( .OUT(na557_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na90_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b1), .IN8(~na1024_1),
                     .CINX(1'b0), .CINY1(na555_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y70     80'h00_0078_00_0020_0C66_C55C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a559_1 ( .OUT(na559_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na720_1), .IN6(1'b1), .IN7(1'b1), .IN8(na925_2),
                     .CINX(1'b0), .CINY1(na582_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a559_4 ( .OUT(na559_2), .COUTY1(na559_4), .IN1(1'b1), .IN2(na889_2), .IN3(~na721_1), .IN4(1'b1), .IN5(~na720_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na925_2), .CINX(1'b0), .CINY1(na582_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y75     80'h00_0078_00_0020_0C66_5C5C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a560_1 ( .OUT(na560_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na935_2), .IN7(~na1714_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na573_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a560_4 ( .OUT(na560_2), .COUTY1(na560_4), .IN1(1'b1), .IN2(na899_2), .IN3(~na731_1), .IN4(1'b1), .IN5(1'b1), .IN6(na935_2),
                     .IN7(~na1714_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na573_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y76     80'h00_0078_00_0020_0C66_3A3C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a562_1 ( .OUT(na562_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na937_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na732_2),
                     .CINX(1'b0), .CINY1(na560_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a562_4 ( .OUT(na562_2), .COUTY1(na562_4), .IN1(1'b1), .IN2(na901_2), .IN3(1'b1), .IN4(~na733_1), .IN5(na937_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(~na732_2), .CINX(1'b0), .CINY1(na560_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y77     80'h00_0078_00_0020_0C66_3AA5
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a564_1 ( .OUT(na564_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na734_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1721_2),
                     .CINX(1'b0), .CINY1(na562_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a564_4 ( .OUT(na564_2), .IN1(~na735_1), .IN2(1'b1), .IN3(na940_2), .IN4(1'b1), .IN5(na734_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na1721_2),
                     .CINX(1'b0), .CINY1(na562_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y71     80'h00_0078_00_0020_0C66_A53C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a567_1 ( .OUT(na567_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na722_2), .IN6(1'b1), .IN7(na927_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na559_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a567_4 ( .OUT(na567_2), .COUTY1(na567_4), .IN1(1'b1), .IN2(na891_2), .IN3(1'b1), .IN4(~na723_1), .IN5(~na722_2), .IN6(1'b1),
                     .IN7(na927_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na559_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y72     80'h00_0078_00_0020_0C66_C53C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a569_1 ( .OUT(na569_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na724_1), .IN6(1'b1), .IN7(1'b1), .IN8(na929_1),
                     .CINX(1'b0), .CINY1(na567_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a569_4 ( .OUT(na569_2), .COUTY1(na569_4), .IN1(1'b1), .IN2(na893_2), .IN3(1'b1), .IN4(~na725_1), .IN5(~na724_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na929_1), .CINX(1'b0), .CINY1(na567_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y73     80'h00_0078_00_0020_0C66_5A3A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a571_1 ( .OUT(na571_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na931_1), .IN6(1'b1), .IN7(~na726_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na569_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a571_4 ( .OUT(na571_2), .COUTY1(na571_4), .IN1(na895_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1710_2), .IN5(na931_1), .IN6(1'b1),
                     .IN7(~na726_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na569_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x51y74     80'h00_0078_00_0020_0C66_C33A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a573_1 ( .OUT(na573_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na728_1), .IN7(1'b1), .IN8(na933_2),
                     .CINX(1'b0), .CINY1(na571_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a573_4 ( .OUT(na573_2), .COUTY1(na573_4), .IN1(na897_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1712_2), .IN5(1'b1), .IN6(~na728_1),
                     .IN7(1'b1), .IN8(na933_2), .CINX(1'b0), .CINY1(na571_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x24y53     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a575_2 ( .OUT(na575_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a575_6 ( .COUTY1(na575_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na575_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x35y74     80'h00_0078_00_0020_0C66_CA05
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a576_1 ( .OUT(na576_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na62_1), .IN6(1'b1), .IN7(1'b1), .IN8(na60_1),
                     .CINX(1'b0), .CINY1(na587_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a576_4 ( .OUT(na576_2), .COUTY1(na576_4), .IN1(~na64_2), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(na62_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na60_1), .CINX(1'b0), .CINY1(na587_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x35y75     80'h00_0078_00_0020_0C66_0C03
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a578_1 ( .OUT(na578_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na66_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na576_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a578_4 ( .OUT(na578_2), .COUTY1(na578_4), .IN1(1'b1), .IN2(~na68_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na66_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na576_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x35y76     80'h00_0018_00_0010_0666_000A
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a580_1 ( .OUT(na580_1), .COUTY1(na580_4), .IN1(na70_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na578_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x51y53     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a581_2 ( .OUT(na581_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a581_6 ( .COUTY1(na581_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na581_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x51y69     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a582_2 ( .OUT(na582_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a582_6 ( .COUTY1(na582_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na582_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x51y48     80'h00_FA60_00_0020_0C66_CCC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a583_1 ( .OUT(na583_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na583_1), .IN7(1'b1), .IN8(na866_2),
                     .CINX(1'b0), .CINY1(na599_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a583_2 ( .OUT(na583_1), .CLK(na624_1), .EN(na169_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na583_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a583_4 ( .OUT(na583_2), .COUTY1(na583_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na866_1), .IN5(1'b1), .IN6(na583_1), .IN7(1'b1),
                     .IN8(na866_2), .CINX(1'b0), .CINY1(na599_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x51y49     80'h00_FA60_00_0020_0C66_0AA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a585_1 ( .OUT(na585_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na585_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na583_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a585_2 ( .OUT(na585_1), .CLK(na624_1), .EN(na169_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na585_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a585_4 ( .OUT(na585_2), .IN1(1'b0), .IN2(1'b0), .IN3(na868_1), .IN4(1'b1), .IN5(na585_1), .IN6(1'b1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na583_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x35y73     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a587_2 ( .OUT(na587_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a587_6 ( .COUTY1(na587_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na587_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF////      x56y58     80'h00_0018_00_0010_0666_000C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a589_1 ( .OUT(na589_1), .IN1(1'b1), .IN2(na82_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na598_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x56y53     80'h00_0078_00_0020_0C66_AC0A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a590_1 ( .OUT(na590_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na876_2), .IN7(na72_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na610_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a590_4 ( .OUT(na590_2), .COUTY1(na590_4), .IN1(na73_1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na876_2), .IN7(na72_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na610_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x56y54     80'h00_0078_00_0020_0C66_FCCF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a592_1 ( .OUT(na592_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na74_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na590_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a592_4 ( .OUT(na592_2), .COUTY1(na592_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na75_1), .IN5(1'b1), .IN6(na74_1), .IN7(1'b1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na590_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x56y55     80'h00_0078_00_0020_0C66_CFC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a594_1 ( .OUT(na594_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na76_1),
                     .CINX(1'b0), .CINY1(na592_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a594_4 ( .OUT(na594_2), .COUTY1(na594_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na77_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na76_1), .CINX(1'b0), .CINY1(na592_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x56y56     80'h00_0078_00_0020_0C66_A00C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a596_1 ( .OUT(na596_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na78_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na594_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a596_4 ( .OUT(na596_2), .COUTY1(na596_4), .IN1(1'b1), .IN2(na79_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na78_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na594_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x56y57     80'h00_0078_00_0020_0C66_0CC0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a598_1 ( .OUT(na598_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na80_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na596_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a598_4 ( .OUT(na598_2), .COUTY1(na598_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(na81_1), .IN5(1'b1), .IN6(na80_1), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na596_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x51y47     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a599_2 ( .OUT(na599_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a599_6 ( .COUTY1(na599_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na599_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x57y53     80'h00_0078_00_0020_0C66_AACF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a601_1 ( .OUT(na601_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1693_2), .IN6(1'b1), .IN7(na590_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na615_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a601_4 ( .OUT(na601_2), .COUTY1(na601_4), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na592_1), .IN5(na1693_2), .IN6(1'b1),
                     .IN7(na590_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na615_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x57y54     80'h00_0078_00_0020_0C66_CFA0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a603_1 ( .OUT(na603_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na592_2),
                     .CINX(1'b0), .CINY1(na601_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a603_4 ( .OUT(na603_2), .COUTY1(na603_4), .IN1(1'b0), .IN2(1'b1), .IN3(na594_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na592_2), .CINX(1'b0), .CINY1(na601_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x57y55     80'h00_0078_00_0020_0C66_A0C0
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a605_1 ( .OUT(na605_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(na594_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na603_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a605_4 ( .OUT(na605_2), .COUTY1(na605_4), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(na596_1), .IN5(1'b0), .IN6(1'b1), .IN7(na594_2),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na603_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x57y56     80'h00_0078_00_0020_0C66_CFAF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a607_1 ( .OUT(na607_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na596_2),
                     .CINX(1'b0), .CINY1(na605_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a607_4 ( .OUT(na607_2), .COUTY1(na607_4), .IN1(1'b1), .IN2(1'b1), .IN3(na598_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na596_2), .CINX(1'b0), .CINY1(na605_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x57y57     80'h00_0078_00_0020_0C66_A0CF
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a609_1 ( .OUT(na609_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b1), .IN7(na598_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na607_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a609_4 ( .OUT(na609_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na589_1), .IN5(1'b0), .IN6(1'b1), .IN7(na598_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na607_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x56y52     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a610_2 ( .OUT(na610_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a610_6 ( .COUTY1(na610_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na610_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2/D//ADDF2/      x29y79     80'h00_FA60_00_0020_0C66_CA0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a611_1 ( .OUT(na611_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na611_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1744_2),
                     .CINX(1'b0), .CINY1(na621_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a611_2 ( .OUT(na611_1), .CLK(na624_1), .EN(na171_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na611_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a611_4 ( .OUT(na611_2), .COUTY1(na611_4), .IN1(1'b1), .IN2(na871_2), .IN3(1'b0), .IN4(1'b0), .IN5(na611_1), .IN6(1'b1), .IN7(1'b1),
                     .IN8(na1744_2), .CINX(1'b0), .CINY1(na621_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x29y80     80'h00_FA60_00_0020_0C66_0C0C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a613_1 ( .OUT(na613_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na613_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na611_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a613_2 ( .OUT(na613_1), .CLK(na624_1), .EN(na171_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na613_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a613_4 ( .OUT(na613_2), .IN1(1'b1), .IN2(na875_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na613_1), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na611_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x57y52     80'h00_3F00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a615_2 ( .OUT(na615_1), .CLK(1'b1), .EN(1'b0), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a615_6 ( .COUTY1(na615_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na615_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x26y73     80'h00_0078_00_0020_0C66_3330
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a616_1 ( .OUT(na616_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na1025_1), .IN7(1'b1), .IN8(~na1026_1),
                     .CINX(1'b0), .CINY1(na941_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a616_4 ( .OUT(na616_2), .COUTY1(na616_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1027_1), .IN5(1'b1), .IN6(~na1025_1),
                     .IN7(1'b1), .IN8(~na1026_1), .CINX(1'b0), .CINY1(na941_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x26y74     80'h00_0078_00_0020_0C66_5050
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a618_1 ( .OUT(na618_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(~na1028_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na616_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a618_4 ( .OUT(na618_2), .COUTY1(na618_4), .IN1(1'b0), .IN2(1'b0), .IN3(~na1029_2), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(~na1028_1),
                     .IN8(1'b1), .CINX(1'b0), .CINY1(na616_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF////      x26y75     80'h00_0018_00_0010_0666_0030
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a620_1 ( .OUT(na620_1), .COUTY1(na620_4), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na1030_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na618_4), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x29y78     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a621_2 ( .OUT(na621_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a621_6 ( .COUTY1(na621_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na621_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
GLBOUT     #(.GLBOUT_CFG (64'h0000_0000_0014_0014)) 
           _a624 ( .GLB0(na624_1), .GLB1(na624_2), .GLB2(_d0), .GLB3(_d1), .CLK_FB0(_d2), .CLK_FB1(_d3), .CLK_FB2(_d4), .CLK_FB3(_d5),
                   .CLK0_0(na1038_6), .CLK0_90(na1038_5), .CLK0_180(na1038_4), .CLK0_270(na1038_3), .CLK0_BYP(1'b0), .CLK1_0(na1039_6),
                   .CLK1_90(na1039_5), .CLK1_180(na1039_4), .CLK1_270(na1039_3), .CLK1_BYP(1'b0), .CLK2_0(1'b0), .CLK2_90(1'b0), .CLK2_180(1'b0),
                   .CLK2_270(1'b0), .CLK2_BYP(1'b0), .CLK3_0(1'b0), .CLK3_90(1'b0), .CLK3_180(1'b0), .CLK3_270(1'b0), .CLK3_BYP(1'b0),
                   .USR_GLB0(1'b0), .USR_GLB1(1'b0), .USR_GLB2(1'b0), .USR_GLB3(1'b0), .USR_FB0(1'b0), .USR_FB1(1'b0), .USR_FB2(1'b0),
                   .USR_FB3(1'b0) );
// C_///AND/D      x39y48     80'h00_FE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a634_4 ( .OUT(na634_2_i), .IN1(1'b1), .IN2(na949_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a634_5 ( .OUT(na634_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na634_2_i) );
// C_AND/D///      x39y48     80'h00_FE00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a635_1 ( .OUT(na635_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na949_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a635_2 ( .OUT(na635_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na635_1_i) );
// C_AND/D///      x40y49     80'h00_FE00_00_0000_0C88_F5FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a636_1 ( .OUT(na636_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na951_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a636_2 ( .OUT(na636_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na636_1_i) );
// C_AND/D///      x38y46     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a638_1 ( .OUT(na638_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na480_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a638_2 ( .OUT(na638_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na638_1_i) );
// C_///AND/D      x38y46     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a640_4 ( .OUT(na640_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na489_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a640_5 ( .OUT(na640_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na640_2_i) );
// C_AND/D///      x38y47     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a642_1 ( .OUT(na642_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na491_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a642_2 ( .OUT(na642_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na642_1_i) );
// C_///AND/D      x38y47     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a644_4 ( .OUT(na644_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na493_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a644_5 ( .OUT(na644_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na644_2_i) );
// C_AND/D///      x40y47     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a646_1 ( .OUT(na646_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na495_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a646_2 ( .OUT(na646_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na646_1_i) );
// C_///AND/D      x40y48     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a648_4 ( .OUT(na648_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na471_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a648_5 ( .OUT(na648_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na648_2_i) );
// C_AND/D///      x42y50     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a650_1 ( .OUT(na650_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na473_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a650_2 ( .OUT(na650_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na650_1_i) );
// C_///AND/D      x40y49     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a652_4 ( .OUT(na652_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na475_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a652_5 ( .OUT(na652_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na652_2_i) );
// C_AND/D///      x42y49     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a654_1 ( .OUT(na654_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na477_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a654_2 ( .OUT(na654_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na654_1_i) );
// C_///AND/D      x42y49     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a656_4 ( .OUT(na656_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na479_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a656_5 ( .OUT(na656_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na656_2_i) );
// C_AND/D///      x45y49     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a658_1 ( .OUT(na658_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na482_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a658_2 ( .OUT(na658_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na658_1_i) );
// C_///AND/D      x45y49     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a660_4 ( .OUT(na660_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na484_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a660_5 ( .OUT(na660_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na660_2_i) );
// C_AND/D///      x28y60     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a662_1 ( .OUT(na662_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na486_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a662_2 ( .OUT(na662_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na662_1_i) );
// C_///AND/D      x45y48     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a663_4 ( .OUT(na663_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na173_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a663_5 ( .OUT(na663_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na663_2_i) );
// C_AND/D//AND/D      x58y61     80'h00_FE00_80_0000_0C88_FC5F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a696_1 ( .OUT(na696_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na503_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a696_2 ( .OUT(na696_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na696_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a696_4 ( .OUT(na696_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na696_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a696_5 ( .OUT(na696_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na696_2_i) );
// C_AND/D///      x58y63     80'h00_FE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a698_1 ( .OUT(na698_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na505_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a698_2 ( .OUT(na698_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na698_1_i) );
// C_///AND/D      x56y64     80'h00_FE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a700_4 ( .OUT(na700_2_i), .IN1(1'b1), .IN2(na507_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a700_5 ( .OUT(na700_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na700_2_i) );
// C_AND/D///      x58y64     80'h00_FE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a702_1 ( .OUT(na702_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na509_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a702_2 ( .OUT(na702_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na702_1_i) );
// C_///AND/D      x58y63     80'h00_FE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a704_4 ( .OUT(na704_2_i), .IN1(1'b1), .IN2(na511_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a704_5 ( .OUT(na704_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na704_2_i) );
// C_AND/D///      x58y67     80'h00_FE00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a706_1 ( .OUT(na706_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na498_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a706_2 ( .OUT(na706_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na706_1_i) );
// C_///AND/D      x58y66     80'h00_FE00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a708_4 ( .OUT(na708_2_i), .IN1(1'b1), .IN2(na500_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a708_5 ( .OUT(na708_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na708_2_i) );
// C_AND/D///      x49y67     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a720_1 ( .OUT(na720_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na973_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a720_2 ( .OUT(na720_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na720_1_i) );
// C_AND/D//AND/D      x52y65     80'h00_FA00_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a721_1 ( .OUT(na721_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na721_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a721_2 ( .OUT(na721_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na721_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a721_4 ( .OUT(na721_2_i), .IN1(1'b1), .IN2(na973_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a721_5 ( .OUT(na721_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na721_2_i) );
// C_///AND/D      x49y63     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a722_4 ( .OUT(na722_2_i), .IN1(na981_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a722_5 ( .OUT(na722_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na722_2_i) );
// C_AND/D//AND/D      x54y66     80'h00_FA00_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a723_1 ( .OUT(na723_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na723_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a723_2 ( .OUT(na723_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na723_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a723_4 ( .OUT(na723_2_i), .IN1(na981_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a723_5 ( .OUT(na723_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na723_2_i) );
// C_AND/D///      x51y65     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a724_1 ( .OUT(na724_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na983_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a724_2 ( .OUT(na724_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na724_1_i) );
// C_AND/D//AND/D      x52y66     80'h00_FA00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a725_1 ( .OUT(na725_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na725_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a725_2 ( .OUT(na725_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na725_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a725_4 ( .OUT(na725_2_i), .IN1(1'b1), .IN2(na983_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a725_5 ( .OUT(na725_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na725_2_i) );
// C_///AND/D      x52y67     80'h00_FA00_80_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a726_4 ( .OUT(na726_2_i), .IN1(na985_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a726_5 ( .OUT(na726_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na726_2_i) );
// C_AND/D//AND/D      x55y64     80'h00_FA00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a727_1 ( .OUT(na727_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na727_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a727_2 ( .OUT(na727_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na727_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a727_4 ( .OUT(na727_2_i), .IN1(na985_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a727_5 ( .OUT(na727_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na727_2_i) );
// C_AND/D///      x49y72     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a728_1 ( .OUT(na728_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na987_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a728_2 ( .OUT(na728_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na728_1_i) );
// C_AND/D//AND/D      x51y68     80'h00_FA00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a729_1 ( .OUT(na729_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na729_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a729_2 ( .OUT(na729_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na729_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a729_4 ( .OUT(na729_2_i), .IN1(1'b1), .IN2(na987_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a729_5 ( .OUT(na729_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na729_2_i) );
// C_AND/D///      x49y71     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a730_1 ( .OUT(na730_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na974_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a730_2 ( .OUT(na730_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na730_1_i) );
// C_AND/D//AND/D      x58y77     80'h00_FA00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a731_1 ( .OUT(na731_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na731_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a731_2 ( .OUT(na731_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na731_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a731_4 ( .OUT(na731_2_i), .IN1(na974_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a731_5 ( .OUT(na731_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na731_2_i) );
// C_///AND/D      x52y78     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a732_4 ( .OUT(na732_2_i), .IN1(1'b1), .IN2(na976_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a732_5 ( .OUT(na732_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na732_2_i) );
// C_AND/D//AND/D      x52y80     80'h00_FA00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a733_1 ( .OUT(na733_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na733_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a733_2 ( .OUT(na733_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na733_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a733_4 ( .OUT(na733_2_i), .IN1(1'b1), .IN2(na976_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a733_5 ( .OUT(na733_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na733_2_i) );
// C_AND/D//AND/D      x51y79     80'h00_FA00_80_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a734_1 ( .OUT(na734_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na978_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a734_2 ( .OUT(na734_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na734_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a734_4 ( .OUT(na734_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na962_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a734_5 ( .OUT(na734_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na734_2_i) );
// C_AND/D///      x45y73     80'h00_FA00_00_0000_0C88_FCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a735_1 ( .OUT(na735_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na979_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a735_2 ( .OUT(na735_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na735_1_i) );
// C_///AND/D      x54y61     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a744_4 ( .OUT(na744_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na434_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a744_5 ( .OUT(na744_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na744_2_i) );
// C_AND/D//AND/D      x49y62     80'h00_FE00_80_0000_0C88_AFF3
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a745_1 ( .OUT(na745_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na434_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a745_2 ( .OUT(na745_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na745_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a745_4 ( .OUT(na745_2_i), .IN1(1'b1), .IN2(~na745_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a745_5 ( .OUT(na745_2), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na745_2_i) );
// C_AND/D///      x54y50     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a748_1 ( .OUT(na748_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na512_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a748_2 ( .OUT(na748_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na748_1_i) );
// C_///AND/D      x54y47     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a750_4 ( .OUT(na750_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na532_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a750_5 ( .OUT(na750_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na750_2_i) );
// C_AND/D///      x58y51     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a752_1 ( .OUT(na752_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na534_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a752_2 ( .OUT(na752_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na752_1_i) );
// C_AND/D///      x56y51     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a754_1 ( .OUT(na754_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na536_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a754_2 ( .OUT(na754_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na754_1_i) );
// C_///AND/D      x54y51     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a756_4 ( .OUT(na756_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na538_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a756_5 ( .OUT(na756_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na756_2_i) );
// C_///AND/D      x54y57     80'h00_FE00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a758_4 ( .OUT(na758_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na513_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a758_5 ( .OUT(na758_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na758_2_i) );
// C_///AND/D      x58y57     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a760_4 ( .OUT(na760_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na515_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a760_5 ( .OUT(na760_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na760_2_i) );
// C_AND/D///      x54y55     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a762_1 ( .OUT(na762_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na517_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a762_2 ( .OUT(na762_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na762_1_i) );
// C_///AND/D      x54y59     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a764_4 ( .OUT(na764_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na519_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a764_5 ( .OUT(na764_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na764_2_i) );
// C_AND/D///      x49y55     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a766_1 ( .OUT(na766_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na521_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a766_2 ( .OUT(na766_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na766_1_i) );
// C_AND/D///      x51y58     80'h00_FE00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a768_1 ( .OUT(na768_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na524_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a768_2 ( .OUT(na768_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na768_1_i) );
// C_AND/D///      x54y59     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a770_1 ( .OUT(na770_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na526_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a770_2 ( .OUT(na770_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na770_1_i) );
// C_///AND/D      x54y62     80'h00_FE00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a772_4 ( .OUT(na772_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na528_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a772_5 ( .OUT(na772_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na772_2_i) );
// C_AND/D///      x57y47     80'h00_FE00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a774_1 ( .OUT(na774_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na530_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a774_2 ( .OUT(na774_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na774_1_i) );
// C_AND/D//AND/D      x44y56     80'h00_FE00_80_0000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a775_1 ( .OUT(na775_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na775_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a775_2 ( .OUT(na775_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na775_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a775_4 ( .OUT(na775_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1482_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a775_5 ( .OUT(na775_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na775_2_i) );
// C_AND/D//AND/D      x49y50     80'h00_FE00_80_0000_0C88_FCCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a776_1 ( .OUT(na776_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na776_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a776_2 ( .OUT(na776_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na776_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a776_4 ( .OUT(na776_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na1482_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a776_5 ( .OUT(na776_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na776_2_i) );
// C_AND/D//AND/D      x44y57     80'h00_FE00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a777_1 ( .OUT(na777_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na777_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a777_2 ( .OUT(na777_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na777_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a777_4 ( .OUT(na777_2_i), .IN1(na1504_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a777_5 ( .OUT(na777_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na777_2_i) );
// C_AND/D//AND/D      x49y54     80'h00_FE00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a778_1 ( .OUT(na778_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na778_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a778_2 ( .OUT(na778_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na778_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a778_4 ( .OUT(na778_2_i), .IN1(na1504_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a778_5 ( .OUT(na778_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na778_2_i) );
// C_AND/D//AND/D      x44y58     80'h00_FE00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a779_1 ( .OUT(na779_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na779_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a779_2 ( .OUT(na779_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na779_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a779_4 ( .OUT(na779_2_i), .IN1(1'b1), .IN2(na1505_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a779_5 ( .OUT(na779_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na779_2_i) );
// C_AND/D//AND/D      x49y57     80'h00_FE00_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a780_1 ( .OUT(na780_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na780_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a780_2 ( .OUT(na780_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na780_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a780_4 ( .OUT(na780_2_i), .IN1(1'b1), .IN2(na1505_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a780_5 ( .OUT(na780_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na780_2_i) );
// C_AND/D//AND/D      x44y59     80'h00_FE00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a781_1 ( .OUT(na781_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na781_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a781_2 ( .OUT(na781_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na781_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a781_4 ( .OUT(na781_2_i), .IN1(na1506_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a781_5 ( .OUT(na781_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na781_2_i) );
// C_AND/D//AND/D      x49y56     80'h00_FE00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a782_1 ( .OUT(na782_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na782_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a782_2 ( .OUT(na782_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na782_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a782_4 ( .OUT(na782_2_i), .IN1(na1506_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a782_5 ( .OUT(na782_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na782_2_i) );
// C_AND/D//AND/D      x44y60     80'h00_FE00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a783_1 ( .OUT(na783_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na783_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a783_2 ( .OUT(na783_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na783_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a783_4 ( .OUT(na783_2_i), .IN1(1'b1), .IN2(na1507_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a783_5 ( .OUT(na783_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na783_2_i) );
// C_AND/D//AND/D      x51y57     80'h00_FE00_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a784_1 ( .OUT(na784_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na784_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a784_2 ( .OUT(na784_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na784_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a784_4 ( .OUT(na784_2_i), .IN1(1'b1), .IN2(na1507_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a784_5 ( .OUT(na784_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na784_2_i) );
// C_AND/D//AND/D      x44y61     80'h00_FE00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a785_1 ( .OUT(na785_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na785_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a785_2 ( .OUT(na785_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na785_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a785_4 ( .OUT(na785_2_i), .IN1(na1508_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a785_5 ( .OUT(na785_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na785_2_i) );
// C_AND/D//AND/D      x53y57     80'h00_FE00_80_0000_0C88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a786_1 ( .OUT(na786_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na786_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a786_2 ( .OUT(na786_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na786_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a786_4 ( .OUT(na786_2_i), .IN1(na1508_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a786_5 ( .OUT(na786_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na786_2_i) );
// C_AND/D//AND/D      x44y62     80'h00_FE00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a787_1 ( .OUT(na787_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na787_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a787_2 ( .OUT(na787_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na787_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a787_4 ( .OUT(na787_2_i), .IN1(1'b1), .IN2(na1509_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a787_5 ( .OUT(na787_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na787_2_i) );
// C_AND/D//AND/D      x49y58     80'h00_FE00_80_0000_0C88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a788_1 ( .OUT(na788_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na788_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a788_2 ( .OUT(na788_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na788_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a788_4 ( .OUT(na788_2_i), .IN1(1'b1), .IN2(na1509_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a788_5 ( .OUT(na788_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na788_2_i) );
// C_AND/D//AND/D      x44y63     80'h00_FE00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a789_1 ( .OUT(na789_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na789_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a789_2 ( .OUT(na789_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na789_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a789_4 ( .OUT(na789_2_i), .IN1(na1510_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a789_5 ( .OUT(na789_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na789_2_i) );
// C_AND/D//AND/D      x49y60     80'h00_FE00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a790_1 ( .OUT(na790_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na790_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a790_2 ( .OUT(na790_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na790_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a790_4 ( .OUT(na790_2_i), .IN1(na1510_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a790_5 ( .OUT(na790_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na790_2_i) );
// C_AND/D//AND/D      x44y64     80'h00_FE00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a791_1 ( .OUT(na791_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na791_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a791_2 ( .OUT(na791_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na791_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a791_4 ( .OUT(na791_2_i), .IN1(1'b1), .IN2(na1511_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a791_5 ( .OUT(na791_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na791_2_i) );
// C_AND/D//AND/D      x51y59     80'h00_FE00_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a792_1 ( .OUT(na792_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na792_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a792_2 ( .OUT(na792_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na792_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a792_4 ( .OUT(na792_2_i), .IN1(1'b1), .IN2(na1511_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a792_5 ( .OUT(na792_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na792_2_i) );
// C_AND/D//AND/D      x44y65     80'h00_FE00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a793_1 ( .OUT(na793_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na793_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a793_2 ( .OUT(na793_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na793_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a793_4 ( .OUT(na793_2_i), .IN1(na1512_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a793_5 ( .OUT(na793_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na793_2_i) );
// C_AND/D//AND/D      x50y62     80'h00_FE00_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a794_1 ( .OUT(na794_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na794_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a794_2 ( .OUT(na794_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na794_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a794_4 ( .OUT(na794_2_i), .IN1(na1512_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a794_5 ( .OUT(na794_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na794_2_i) );
// C_AND/D//AND/D      x44y66     80'h00_FE00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a795_1 ( .OUT(na795_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na795_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a795_2 ( .OUT(na795_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na795_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a795_4 ( .OUT(na795_2_i), .IN1(1'b1), .IN2(na1513_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a795_5 ( .OUT(na795_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na795_2_i) );
// C_AND/D//AND/D      x50y61     80'h00_FE00_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a796_1 ( .OUT(na796_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na796_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a796_2 ( .OUT(na796_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na796_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a796_4 ( .OUT(na796_2_i), .IN1(1'b1), .IN2(na1513_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a796_5 ( .OUT(na796_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na796_2_i) );
// C_AND/D//AND/D      x44y67     80'h00_FE00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a797_1 ( .OUT(na797_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na797_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a797_2 ( .OUT(na797_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na797_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a797_4 ( .OUT(na797_2_i), .IN1(na1514_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a797_5 ( .OUT(na797_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na797_2_i) );
// C_AND/D//AND/D      x51y62     80'h00_FE00_80_0000_0C88_FCFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a798_1 ( .OUT(na798_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na798_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a798_2 ( .OUT(na798_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na798_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a798_4 ( .OUT(na798_2_i), .IN1(na1514_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a798_5 ( .OUT(na798_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na798_2_i) );
// C_AND/D//AND/D      x44y68     80'h00_FE00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a799_1 ( .OUT(na799_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na799_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a799_2 ( .OUT(na799_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na799_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a799_4 ( .OUT(na799_2_i), .IN1(1'b1), .IN2(na1515_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a799_5 ( .OUT(na799_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na799_2_i) );
// C_AND/D//AND/D      x49y59     80'h00_FE00_80_0000_0C88_FAFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a800_1 ( .OUT(na800_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na800_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a800_2 ( .OUT(na800_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na800_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a800_4 ( .OUT(na800_2_i), .IN1(1'b1), .IN2(na1515_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a800_5 ( .OUT(na800_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na800_2_i) );
// C_AND/D//AND/D      x44y69     80'h00_FE00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a801_1 ( .OUT(na801_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na801_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a801_2 ( .OUT(na801_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na801_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a801_4 ( .OUT(na801_2_i), .IN1(na1516_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a801_5 ( .OUT(na801_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na801_2_i) );
// C_AND/D//AND/D      x50y63     80'h00_FE00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a802_1 ( .OUT(na802_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na802_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a802_2 ( .OUT(na802_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na802_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a802_4 ( .OUT(na802_2_i), .IN1(na1516_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a802_5 ( .OUT(na802_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na802_2_i) );
// C_///AND/D      x33y68     80'h00_FA00_80_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a844_4 ( .OUT(na844_2_i), .IN1(1'b1), .IN2(~na844_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a844_5 ( .OUT(na844_2), .CLK(na624_1), .EN(na156_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na844_2_i) );
// C_AND/D//AND/D      x22y68     80'h00_FA00_80_0000_0C88_AF3F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a862_1 ( .OUT(na862_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na426_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a862_2 ( .OUT(na862_1), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na862_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a862_4 ( .OUT(na862_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na862_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a862_5 ( .OUT(na862_2), .CLK(na624_1), .EN(na168_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na862_2_i) );
// C_AND/D//AND/D      x50y48     80'h00_FA00_80_0000_0C88_FC3F
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a866_1 ( .OUT(na866_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na583_2), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a866_2 ( .OUT(na866_1), .CLK(na624_1), .EN(na169_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na866_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a866_4 ( .OUT(na866_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na866_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a866_5 ( .OUT(na866_2), .CLK(na624_1), .EN(na169_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na866_2_i) );
// C_AND/D///      x50y57     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a868_1 ( .OUT(na868_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na585_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a868_2 ( .OUT(na868_1), .CLK(na624_1), .EN(na169_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na868_1_i) );
// C_AND/D//AND/D      x31y76     80'h00_FA00_80_0000_0C88_F3FA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a871_1 ( .OUT(na871_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na871_1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a871_2 ( .OUT(na871_1), .CLK(na624_1), .EN(na171_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na871_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a871_4 ( .OUT(na871_2_i), .IN1(na611_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a871_5 ( .OUT(na871_2), .CLK(na624_1), .EN(na171_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na871_2_i) );
// C_///AND/D      x33y74     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a875_4 ( .OUT(na875_2_i), .IN1(1'b1), .IN2(na613_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a875_5 ( .OUT(na875_2), .CLK(na624_1), .EN(na171_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na875_2_i) );
// C_///AND/D      x55y54     80'h00_FD00_80_0000_0C08_FFF3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a876_4 ( .OUT(na876_2_i), .IN1(1'b1), .IN2(~na876_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a876_5 ( .OUT(na876_2), .CLK(~na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na876_2_i) );
// C_AND/D//AND/D      x59y68     80'h00_FA00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a889_1 ( .OUT(na889_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na957_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a889_2 ( .OUT(na889_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na889_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a889_4 ( .OUT(na889_2_i), .IN1(1'b1), .IN2(na889_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a889_5 ( .OUT(na889_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na889_2_i) );
// C_AND/D//AND/D      x51y66     80'h00_FA00_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a891_1 ( .OUT(na891_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na965_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a891_2 ( .OUT(na891_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na891_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a891_4 ( .OUT(na891_2_i), .IN1(1'b1), .IN2(na891_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a891_5 ( .OUT(na891_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na891_2_i) );
// C_AND/D//AND/D      x47y68     80'h00_FA00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a893_1 ( .OUT(na893_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na967_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a893_2 ( .OUT(na893_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na893_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a893_4 ( .OUT(na893_2_i), .IN1(1'b1), .IN2(na893_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a893_5 ( .OUT(na893_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na893_2_i) );
// C_AND/D//AND/D      x47y69     80'h00_FA00_80_0000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a895_1 ( .OUT(na895_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na969_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a895_2 ( .OUT(na895_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na895_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a895_4 ( .OUT(na895_2_i), .IN1(na895_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a895_5 ( .OUT(na895_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na895_2_i) );
// C_AND/D//AND/D      x49y69     80'h00_FA00_80_0000_0C88_CFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a897_1 ( .OUT(na897_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na971_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a897_2 ( .OUT(na897_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na897_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a897_4 ( .OUT(na897_2_i), .IN1(na897_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a897_5 ( .OUT(na897_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na897_2_i) );
// C_AND/D//AND/D      x51y82     80'h00_FA00_80_0000_0C88_AFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a899_1 ( .OUT(na899_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na958_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a899_2 ( .OUT(na899_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na899_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a899_4 ( .OUT(na899_2_i), .IN1(1'b1), .IN2(na899_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a899_5 ( .OUT(na899_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na899_2_i) );
// C_AND/D//AND/D      x53y80     80'h00_FA00_80_0000_0C88_CFFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a901_1 ( .OUT(na901_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na960_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a901_2 ( .OUT(na901_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na901_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a901_4 ( .OUT(na901_2_i), .IN1(1'b1), .IN2(na901_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a901_5 ( .OUT(na901_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na901_2_i) );
// C_///AND/D      x44y53     80'h00_FA00_80_0000_0C08_FF5F
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a904_4 ( .OUT(na904_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(~na904_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0100)) 
           _a904_5 ( .OUT(na904_2), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na904_2_i) );
// C_///AND/D      x44y55     80'h00_FA00_80_0000_0C08_FFFC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a906_4 ( .OUT(na906_2_i), .IN1(1'b1), .IN2(na429_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b1_0000_0100)) 
           _a906_5 ( .OUT(na906_2), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na906_2_i) );
// C_AND/D///      x45y55     80'h00_FA00_00_0000_0C88_FAFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a908_1 ( .OUT(na908_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na431_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'b0_0000_0000)) 
           _a908_2 ( .OUT(na908_1), .CLK(na624_1), .EN(na82_1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na908_1_i) );
// C_///AND/D      x54y68     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a925_4 ( .OUT(na925_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na957_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a925_5 ( .OUT(na925_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na925_2_i) );
// C_///AND/D      x52y69     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a927_4 ( .OUT(na927_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na965_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a927_5 ( .OUT(na927_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na927_2_i) );
// C_AND/D///      x52y70     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a929_1 ( .OUT(na929_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na967_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a929_2 ( .OUT(na929_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na929_1_i) );
// C_AND/D///      x41y75     80'h00_FA00_00_0000_0C88_AFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a931_1 ( .OUT(na931_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na969_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a931_2 ( .OUT(na931_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na931_1_i) );
// C_///AND/D      x42y78     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a933_4 ( .OUT(na933_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na971_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a933_5 ( .OUT(na933_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na933_2_i) );
// C_///AND/D      x43y78     80'h00_FA00_80_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a935_4 ( .OUT(na935_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na958_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a935_5 ( .OUT(na935_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na935_2_i) );
// C_AND/D///      x55y79     80'h00_FA00_00_0000_0C88_CFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a937_1 ( .OUT(na937_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na960_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a937_2 ( .OUT(na937_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na937_1_i) );
// C_///AND/D      x56y81     80'h00_FA00_80_0000_0C08_FFCF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a940_4 ( .OUT(na940_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na963_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a940_5 ( .OUT(na940_2), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na940_2_i) );
// C_/C_0_1///      x26y72     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a941_2 ( .OUT(na941_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a941_6 ( .COUTY1(na941_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na941_1),
                     .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_ADDF2///ADDF2/      x47y60     80'h00_0078_00_0020_0C66_AACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a942_1 ( .OUT(na942_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na256_2), .IN6(1'b1), .IN7(na202_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na955_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a942_4 ( .OUT(na942_2), .COUTY1(na942_4), .IN1(na256_1), .IN2(1'b1), .IN3(1'b1), .IN4(na211_1), .IN5(na256_2), .IN6(1'b1),
                     .IN7(na202_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na955_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x47y61     80'h00_0078_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a944_1 ( .OUT(na944_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na258_2), .IN6(1'b1), .IN7(na220_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na942_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a944_4 ( .OUT(na944_2), .COUTY1(na944_4), .IN1(na258_1), .IN2(1'b1), .IN3(na229_1), .IN4(1'b1), .IN5(na258_2), .IN6(1'b1),
                     .IN7(na220_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na942_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x47y62     80'h00_0078_00_0020_0C66_ACAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a946_1 ( .OUT(na946_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na259_2), .IN7(na238_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na944_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a946_4 ( .OUT(na946_2), .IN1(na260_1), .IN2(1'b1), .IN3(na244_1), .IN4(1'b1), .IN5(1'b1), .IN6(na259_2), .IN7(na238_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na944_4), .PINX(1'b0), .PINY1(1'b0) );
// C_C_XOR////      x45y70     80'h00_0018_00_0010_0666_0006
C_C_XOR    #(.CPE_CFG (9'b0_0010_0000)) 
           _a948_1 ( .OUT(na948_1), .IN1(na415_1), .IN2(na414_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na415_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x47y56     80'h00_0078_00_0020_0C66_4A4A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a949_1 ( .OUT(na949_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na290_2), .IN6(1'b1), .IN7(~na177_1), .IN8(na1092_2),
                     .CINX(1'b0), .CINY1(na1036_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a949_4 ( .OUT(na949_2), .COUTY1(na949_4), .IN1(na290_1), .IN2(1'b1), .IN3(~na267_1), .IN4(na1092_1), .IN5(na290_2), .IN6(1'b1),
                     .IN7(~na177_1), .IN8(na1092_2), .CINX(1'b0), .CINY1(na1036_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x47y57     80'h00_0078_00_0020_0C66_C24A
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a951_1 ( .OUT(na951_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1095_2), .IN6(~na272_1), .IN7(1'b1), .IN8(na292_2),
                     .CINX(1'b0), .CINY1(na949_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a951_4 ( .OUT(na951_2), .COUTY1(na951_4), .IN1(na1671_2), .IN2(1'b1), .IN3(~na1669_2), .IN4(na1805_2), .IN5(na1095_2), .IN6(~na272_1),
                     .IN7(1'b1), .IN8(na292_2), .CINX(1'b0), .CINY1(na949_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x47y58     80'h00_0078_00_0020_0C66_A44C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a953_1 ( .OUT(na953_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(~na282_1), .IN6(na252_2), .IN7(na293_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na951_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a953_4 ( .OUT(na953_2), .COUTY1(na953_4), .IN1(1'b1), .IN2(na252_1), .IN3(~na288_1), .IN4(na1097_1), .IN5(~na282_1), .IN6(na252_2),
                     .IN7(na293_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na951_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2///ADDF2/      x47y59     80'h00_0078_00_0020_0C66_CAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a955_1 ( .OUT(na955_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na254_2), .IN6(1'b1), .IN7(1'b1), .IN8(na178_1),
                     .CINX(1'b0), .CINY1(na953_4), .PINX(1'b0), .PINY1(1'b0) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a955_4 ( .OUT(na955_2), .COUTY1(na955_4), .IN1(na254_1), .IN2(1'b1), .IN3(na193_1), .IN4(1'b1), .IN5(na254_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na178_1), .CINX(1'b0), .CINY1(na953_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x54y70     80'h00_FA60_00_0020_0C66_A3CA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a957_1 ( .OUT(na957_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(~na893_1), .IN7(na319_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na1037_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a957_2 ( .OUT(na957_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na957_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a957_4 ( .OUT(na957_2), .COUTY1(na957_4), .IN1(na120_1), .IN2(1'b1), .IN3(1'b1), .IN4(na300_1), .IN5(1'b1), .IN6(~na893_1),
                     .IN7(na319_1), .IN8(1'b1), .CINX(1'b0), .CINY1(na1037_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x54y75     80'h00_FA60_00_0020_0C66_AAC2
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a958_1 ( .OUT(na958_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1098_2), .IN6(1'b1), .IN7(na312_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na971_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a958_2 ( .OUT(na958_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na958_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a958_4 ( .OUT(na958_2), .COUTY1(na958_4), .IN1(na1098_1), .IN2(~na295_1), .IN3(1'b1), .IN4(na314_1), .IN5(na1098_2), .IN6(1'b1),
                     .IN7(na312_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na971_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x/D//ADDF2x/      x54y76     80'h00_FA60_00_0020_0C66_9AA9
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a960_1 ( .OUT(na960_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na296_1), .IN6(1'b0), .IN7(na1112_2), .IN8(~na960_1),
                     .CINX(1'b0), .CINY1(na958_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a960_2 ( .OUT(na960_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na960_1_i) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a960_4 ( .OUT(na960_2), .COUTY1(na960_4), .IN1(na1806_2), .IN2(~na901_1), .IN3(na297_1), .IN4(1'b0), .IN5(na296_1), .IN6(1'b0),
                     .IN7(na1112_2), .IN8(~na960_1), .CINX(1'b0), .CINY1(na958_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDFx/D///      x54y77     80'h00_FA00_00_0010_0666_009A
C_ADDFx    #(.CPE_CFG (9'b0_0010_0000)) 
           _a962_1 ( .OUT(na962_1_i), .COUTY1(na962_4), .IN1(na298_1), .IN2(1'b0), .IN3(~na962_1), .IN4(na1113_2), .IN5(1'b0), .IN6(1'b0),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na960_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a962_2 ( .OUT(na962_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na962_1_i) );
// C_ADDF/D///      x54y78     80'h00_FA00_00_0010_0666_005C
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a963_1 ( .OUT(na963_1_i), .IN1(1'b1), .IN2(na299_1), .IN3(~na318_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na962_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a963_2 ( .OUT(na963_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na963_1_i) );
// C_ADDF2/D//ADDF2/      x54y71     80'h00_FA60_00_0020_0C66_5ACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a965_1 ( .OUT(na965_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na122_1), .IN6(1'b1), .IN7(~na304_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na957_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a965_2 ( .OUT(na965_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na965_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a965_4 ( .OUT(na965_2), .COUTY1(na965_4), .IN1(na124_2), .IN2(1'b1), .IN3(1'b1), .IN4(na305_1), .IN5(na122_1), .IN6(1'b1),
                     .IN7(~na304_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na957_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x54y72     80'h00_FA60_00_0020_0C66_CCCC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a967_1 ( .OUT(na967_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na307_2), .IN7(1'b1), .IN8(na128_2),
                     .CINX(1'b0), .CINY1(na965_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a967_2 ( .OUT(na967_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na967_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a967_4 ( .OUT(na967_2), .COUTY1(na967_4), .IN1(1'b1), .IN2(na307_1), .IN3(1'b1), .IN4(na128_1), .IN5(1'b1), .IN6(na307_2),
                     .IN7(1'b1), .IN8(na128_2), .CINX(1'b0), .CINY1(na965_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x54y73     80'h00_FA60_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a969_1 ( .OUT(na969_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na132_2), .IN6(1'b1), .IN7(na309_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na967_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a969_2 ( .OUT(na969_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na969_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a969_4 ( .OUT(na969_2), .COUTY1(na969_4), .IN1(na132_1), .IN2(1'b1), .IN3(na309_1), .IN4(1'b1), .IN5(na132_2), .IN6(1'b1),
                     .IN7(na309_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na967_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x54y74     80'h00_FA60_00_0020_0C66_CCCC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a971_1 ( .OUT(na971_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b1), .IN6(na136_2), .IN7(1'b1), .IN8(na311_2),
                     .CINX(1'b0), .CINY1(na969_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a971_2 ( .OUT(na971_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na971_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a971_4 ( .OUT(na971_2), .COUTY1(na971_4), .IN1(1'b1), .IN2(na136_1), .IN3(1'b1), .IN4(na311_1), .IN5(1'b1), .IN6(na136_2),
                     .IN7(1'b1), .IN8(na311_2), .CINX(1'b0), .CINY1(na969_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x53y68     80'h00_FA60_00_0020_0C66_3AAC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a973_1 ( .OUT(na973_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na345_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na725_2),
                     .CINX(1'b0), .CINY1(na1050_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a973_2 ( .OUT(na973_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na973_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a973_4 ( .OUT(na973_2), .COUTY1(na973_4), .IN1(1'b1), .IN2(na138_1), .IN3(na326_1), .IN4(1'b1), .IN5(na345_1), .IN6(1'b1),
                     .IN7(1'b1), .IN8(~na725_2), .CINX(1'b0), .CINY1(na1050_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x53y73     80'h00_FA60_00_0020_0C66_AA2C
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a974_1 ( .OUT(na974_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1114_2), .IN6(1'b1), .IN7(na338_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na987_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a974_2 ( .OUT(na974_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na974_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a974_4 ( .OUT(na974_2), .COUTY1(na974_4), .IN1(1'b1), .IN2(na340_1), .IN3(na1807_2), .IN4(~na321_1), .IN5(na1114_2), .IN6(1'b1),
                     .IN7(na338_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na987_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2x/D//ADDF2x/      x53y74     80'h00_FA60_00_0020_0C66_A99C
C_ADDF2x   #(.CPE_CFG (9'b0_0010_0000)) 
           _a976_1 ( .OUT(na976_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1128_2), .IN6(~na976_1), .IN7(na322_2),
                     .IN8(1'b0), .CINX(1'b0), .CINY1(na974_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a976_2 ( .OUT(na976_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na976_1_i) );
C_ADDF2x   #(.CPE_CFG (9'b0_1000_0000)) 
           _a976_4 ( .OUT(na976_2), .COUTY1(na976_4), .IN1(1'b0), .IN2(na323_1), .IN3(na1808_2), .IN4(~na733_2), .IN5(na1128_2), .IN6(~na976_1),
                     .IN7(na322_2), .IN8(1'b0), .CINX(1'b0), .CINY1(na974_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDFx/D///      x53y75     80'h00_FA00_00_0010_0666_00A9
C_ADDFx    #(.CPE_CFG (9'b0_0010_0000)) 
           _a978_1 ( .OUT(na978_1_i), .COUTY1(na978_4), .IN1(~na978_1), .IN2(na1129_1), .IN3(na324_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0),
                     .IN7(1'b0), .IN8(1'b0), .CINX(1'b0), .CINY1(na976_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a978_2 ( .OUT(na978_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na978_1_i) );
// C_ADDF/D///      x53y76     80'h00_FA00_00_0010_0666_00A3
C_ADDF     #(.CPE_CFG (9'b0_0010_0000)) 
           _a979_1 ( .OUT(na979_1_i), .IN1(1'b1), .IN2(~na344_1), .IN3(na325_1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                     .CINX(1'b0), .CINY1(na978_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a979_2 ( .OUT(na979_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na979_1_i) );
// C_ADDF2/D//ADDF2/      x53y69     80'h00_FA60_00_0020_0C66_5ACC
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a981_1 ( .OUT(na981_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na140_1), .IN6(1'b1), .IN7(~na330_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na973_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a981_2 ( .OUT(na981_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na981_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a981_4 ( .OUT(na981_2), .COUTY1(na981_4), .IN1(1'b1), .IN2(na331_1), .IN3(1'b1), .IN4(na142_1), .IN5(na140_1), .IN6(1'b1),
                     .IN7(~na330_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na973_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x53y70     80'h00_FA60_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a983_1 ( .OUT(na983_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na146_2), .IN6(1'b1), .IN7(na333_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na981_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a983_2 ( .OUT(na983_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na983_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a983_4 ( .OUT(na983_2), .COUTY1(na983_4), .IN1(na146_1), .IN2(1'b1), .IN3(na333_1), .IN4(1'b1), .IN5(na146_2), .IN6(1'b1),
                     .IN7(na333_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na981_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x53y71     80'h00_FA60_00_0020_0C66_CACA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a985_1 ( .OUT(na985_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na335_2), .IN6(1'b1), .IN7(1'b1), .IN8(na150_2),
                     .CINX(1'b0), .CINY1(na983_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a985_2 ( .OUT(na985_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na985_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a985_4 ( .OUT(na985_2), .COUTY1(na985_4), .IN1(na335_1), .IN2(1'b1), .IN3(1'b1), .IN4(na150_1), .IN5(na335_2), .IN6(1'b1),
                     .IN7(1'b1), .IN8(na150_2), .CINX(1'b0), .CINY1(na983_4), .PINX(1'b0), .PINY1(1'b0) );
// C_ADDF2/D//ADDF2/      x53y72     80'h00_FA60_00_0020_0C66_AAAA
C_ADDF2    #(.CPE_CFG (9'b0_0010_0000)) 
           _a987_1 ( .OUT(na987_1_i), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na154_2), .IN6(1'b1), .IN7(na337_2), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(na985_4), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a987_2 ( .OUT(na987_1), .CLK(na624_1), .EN(na172_2), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na987_1_i) );
C_ADDF2    #(.CPE_CFG (9'b0_1000_0000)) 
           _a987_4 ( .OUT(na987_2), .COUTY1(na987_4), .IN1(na154_1), .IN2(1'b1), .IN3(na337_1), .IN4(1'b1), .IN5(na154_2), .IN6(1'b1),
                     .IN7(na337_2), .IN8(1'b1), .CINX(1'b0), .CINY1(na985_4), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x23y81     80'h00_0018_00_0040_0AF3_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a989_1 ( .OUT(na989_1), .IN1(1'b1), .IN2(na98_1), .IN3(1'b1), .IN4(na99_1), .IN5(~na1645_2), .IN6(~na98_2), .IN7(na1641_2),
                     .IN8(na99_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x22y81     80'h00_FE00_00_0040_0AF0_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a990_1 ( .OUT(na990_1_i), .IN1(~na97_1), .IN2(1'b1), .IN3(1'b1), .IN4(na94_2), .IN5(na989_1), .IN6(na9_1), .IN7(na8_1), .IN8(na10_1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a990_2 ( .OUT(na990_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na990_1_i) );
// C_MX4b////      x28y79     80'h00_0018_00_0040_0AF6_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a991_1 ( .OUT(na991_1), .IN1(1'b1), .IN2(~na98_1), .IN3(1'b1), .IN4(na99_1), .IN5(na6_1), .IN6(~na98_2), .IN7(~na8_1), .IN8(na1606_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x19y75     80'h00_0018_00_0040_0AFC_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a992_1 ( .OUT(na992_1), .IN1(1'b1), .IN2(~na98_1), .IN3(1'b1), .IN4(na99_1), .IN5(na6_1), .IN6(na7_2), .IN7(~na4_1), .IN8(~na1612_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x25y74     80'h00_FE00_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a993_1 ( .OUT(na993_1_i), .IN1(na97_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na94_2), .IN5(na992_1), .IN6(na7_2), .IN7(na991_1),
                     .IN8(na11_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a993_2 ( .OUT(na993_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na993_1_i) );
// C_MX4b////      x22y75     80'h00_0018_00_0040_0AF1_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a994_1 ( .OUT(na994_1), .IN1(1'b1), .IN2(na98_1), .IN3(1'b1), .IN4(~na99_1), .IN5(~na6_1), .IN6(na7_2), .IN7(na5_2), .IN8(na1615_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x23y79     80'h00_0018_00_0040_0AFA_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a995_1 ( .OUT(na995_1), .IN1(1'b1), .IN2(~na98_1), .IN3(1'b1), .IN4(na99_1), .IN5(na6_1), .IN6(~na7_2), .IN7(na4_1), .IN8(~na99_2),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x28y74     80'h00_FE00_00_0040_0AF2_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a996_1 ( .OUT(na996_1_i), .IN1(na97_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na94_2), .IN5(na995_1), .IN6(~na98_2), .IN7(na994_1),
                     .IN8(na12_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a996_2 ( .OUT(na996_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na996_1_i) );
// C_MX4b////      x28y80     80'h00_0018_00_0040_0A79_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a997_1 ( .OUT(na997_1), .IN1(1'b1), .IN2(~na98_1), .IN3(1'b1), .IN4(na99_1), .IN5(~na6_1), .IN6(na1614_2), .IN7(na8_1), .IN8(1'b1),
                     .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x25y71     80'h00_FE00_00_0040_0AF2_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a998_1 ( .OUT(na998_1_i), .IN1(na97_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na94_2), .IN5(na14_1), .IN6(~na98_2), .IN7(na13_1),
                     .IN8(na997_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a998_2 ( .OUT(na998_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na998_1_i) );
// C_MX4b////      x20y75     80'h00_0018_00_0040_0AFA_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a999_1 ( .OUT(na999_1), .IN1(1'b1), .IN2(na98_1), .IN3(1'b1), .IN4(na99_1), .IN5(na1607_2), .IN6(~na1610_2), .IN7(na8_1),
                     .IN8(~na99_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x20y78     80'h00_0018_00_0040_0AF9_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1000_1 ( .OUT(na1000_1), .IN1(1'b1), .IN2(~na98_1), .IN3(1'b1), .IN4(na99_1), .IN5(~na1605_2), .IN6(na98_2), .IN7(na8_1),
                      .IN8(~na1642_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x23y74     80'h00_FE00_00_0040_0AF0_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1001_1 ( .OUT(na1001_1_i), .IN1(na97_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na94_2), .IN5(na15_1), .IN6(na98_2), .IN7(na999_1),
                      .IN8(na1000_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1001_2 ( .OUT(na1001_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1001_1_i) );
// C_MX4b////      x23y73     80'h00_0018_00_0040_0AF1_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1002_1 ( .OUT(na1002_1), .IN1(1'b1), .IN2(~na98_1), .IN3(1'b1), .IN4(~na99_1), .IN5(~na1607_2), .IN6(na1608_2), .IN7(na5_2),
                      .IN8(na1606_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x26y77     80'h00_0018_00_0040_0AB2_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1003_1 ( .OUT(na1003_1), .IN1(1'b1), .IN2(na98_1), .IN3(1'b1), .IN4(na99_1), .IN5(na6_1), .IN6(~na98_2), .IN7(1'b0), .IN8(na1609_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x25y75     80'h00_FE00_00_0040_0A70_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1004_1 ( .OUT(na1004_1_i), .IN1(na97_1), .IN2(1'b1), .IN3(1'b1), .IN4(na94_2), .IN5(na1002_1), .IN6(na16_1), .IN7(na1003_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1004_2 ( .OUT(na1004_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1004_1_i) );
// C_MX4b////      x24y74     80'h00_0018_00_0040_0A77_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1005_1 ( .OUT(na1005_1), .IN1(1'b1), .IN2(~na98_1), .IN3(1'b1), .IN4(na99_1), .IN5(~na1645_2), .IN6(~na98_2), .IN7(~na8_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x27y74     80'h00_0018_00_0040_0A7E_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1006_1 ( .OUT(na1006_1), .IN1(1'b1), .IN2(~na98_1), .IN3(1'b1), .IN4(na99_1), .IN5(na6_1), .IN6(~na1610_2), .IN7(~na5_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x27y73     80'h00_FE00_00_0040_0AE1_0035
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1007_1 ( .OUT(na1007_1_i), .IN1(~na97_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na94_2), .IN5(1'b1), .IN6(na1006_1), .IN7(na17_1),
                      .IN8(na1005_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1007_2 ( .OUT(na1007_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1007_1_i) );
// C_MX4b////      x25y78     80'h00_0018_00_0040_0AB6_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1008_1 ( .OUT(na1008_1), .IN1(1'b1), .IN2(~na98_1), .IN3(1'b1), .IN4(na99_1), .IN5(na6_1), .IN6(~na1614_2), .IN7(1'b1), .IN8(na1613_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b/D///      x28y72     80'h00_FE00_00_0040_0AF4_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1009_1 ( .OUT(na1009_1_i), .IN1(~na97_1), .IN2(1'b1), .IN3(1'b1), .IN4(na94_2), .IN5(na18_1), .IN6(na1008_1), .IN7(~na8_1),
                      .IN8(na19_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1009_2 ( .OUT(na1009_1), .CLK(na624_1), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1009_1_i) );
// C_MX4b////      x47y52     80'h00_0018_00_0040_0AF2_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1010_1 ( .OUT(na1010_1), .IN1(~na585_1), .IN2(1'b1), .IN3(~na50_2), .IN4(1'b1), .IN5(na31_2), .IN6(~na51_1), .IN7(na1625_2),
                      .IN8(na1637_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y48     80'h00_0018_00_0040_0AF7_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1011_1 ( .OUT(na1011_1), .IN1(na585_1), .IN2(1'b1), .IN3(1'b1), .IN4(na866_1), .IN5(~na1623_2), .IN6(~na583_1), .IN7(~na26_2),
                      .IN8(na1622_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x45y50     80'h00_0018_00_0040_0AFC_0055
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1012_1 ( .OUT(na1012_1), .IN1(~na585_1), .IN2(1'b1), .IN3(~na50_2), .IN4(1'b1), .IN5(na29_2), .IN6(na53_1), .IN7(~na32_1),
                      .IN8(~na52_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x48y46     80'h00_0018_00_0040_0CE3_3500
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1013_1 ( .OUT(na1013_1), .IN1(na1618_2), .IN2(~na583_1), .IN3(1'b1), .IN4(1'b1), .IN5(~na585_1), .IN6(1'b1), .IN7(1'b1),
                      .IN8(~na866_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x48y49     80'h00_0018_00_0040_0AF0_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1014_1 ( .OUT(na1014_1), .IN1(na585_1), .IN2(1'b1), .IN3(1'b1), .IN4(na866_1), .IN5(na1618_2), .IN6(na25_1), .IN7(na26_2),
                      .IN8(na27_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x49y51     80'h00_0018_00_0040_0AF5_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1015_1 ( .OUT(na1015_1), .IN1(na1739_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1692_2), .IN5(~na1618_2), .IN6(na583_1), .IN7(~na1691_2),
                      .IN8(na866_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y54     80'h00_0018_00_0040_0AFA_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1016_1 ( .OUT(na1016_1), .IN1(na1619_2), .IN2(1'b1), .IN3(~na32_2), .IN4(1'b1), .IN5(na1015_1), .IN6(~na1626_2), .IN7(na1014_1),
                      .IN8(~na24_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x49y49     80'h00_0018_00_0040_0AFB_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1017_1 ( .OUT(na1017_1), .IN1(na1739_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1692_2), .IN5(~na1623_2), .IN6(~na583_1), .IN7(na1691_2),
                      .IN8(~na24_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y52     80'h00_0018_00_0040_0AFB_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1018_1 ( .OUT(na1018_1), .IN1(na585_1), .IN2(1'b1), .IN3(1'b1), .IN4(~na866_1), .IN5(~na1621_2), .IN6(~na583_1), .IN7(na1617_2),
                      .IN8(~na1620_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x49y52     80'h00_0018_00_0040_0AF0_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1019_1 ( .OUT(na1019_1), .IN1(1'b1), .IN2(na1627_2), .IN3(1'b1), .IN4(na24_2), .IN5(na1017_1), .IN6(na1018_1), .IN7(na54_1),
                      .IN8(na28_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_ICOMP////      x50y51     80'h00_0018_00_0000_0C88_C9FF
C_ICOMP    #(.CPE_CFG (9'b0_0000_0000)) 
           _a1020_1 ( .OUT(na1020_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na585_1), .IN6(na1740_2), .IN7(1'b1), .IN8(na23_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x51y51     80'h00_0018_00_0040_0A6B_003A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1021_1 ( .OUT(na1021_1), .IN1(na1739_2), .IN2(1'b1), .IN3(1'b1), .IN4(~na1692_2), .IN5(1'b1), .IN6(~na1616_2), .IN7(na26_2),
                      .IN8(1'b1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y55     80'h00_0018_00_0040_0AF0_005A
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1022_1 ( .OUT(na1022_1), .IN1(na1619_2), .IN2(1'b1), .IN3(~na32_2), .IN4(1'b1), .IN5(na1021_1), .IN6(na1624_2), .IN7(na1020_1),
                      .IN8(na28_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x47y49     80'h00_0018_00_0040_0A66_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1023_1 ( .OUT(na1023_1), .IN1(~na1739_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1692_2), .IN5(1'b0), .IN6(~na25_1), .IN7(~na26_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y56     80'h00_0018_00_0040_0AFC_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1024_1 ( .OUT(na1024_1), .IN1(1'b1), .IN2(na1627_2), .IN3(1'b1), .IN4(na24_2), .IN5(na1023_1), .IN6(na55_1), .IN7(~na56_1),
                      .IN8(~na30_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x37y74     80'h00_0018_00_0040_0A66_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1025_1 ( .OUT(na1025_1), .IN1(1'b1), .IN2(~na871_2), .IN3(1'b1), .IN4(~na1703_2), .IN5(1'b0), .IN6(~na20_2), .IN7(~na21_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x30y76     80'h00_0018_00_0040_0AFD_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1026_1 ( .OUT(na1026_1), .IN1(1'b1), .IN2(~na871_2), .IN3(1'b1), .IN4(~na1703_2), .IN5(~na57_1), .IN6(na871_1), .IN7(~na1743_2),
                      .IN8(~na58_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x30y74     80'h00_0018_00_0040_0AF0_003C
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1027_1 ( .OUT(na1027_1), .IN1(1'b1), .IN2(na613_1), .IN3(1'b1), .IN4(~na1746_2), .IN5(na57_1), .IN6(na20_2), .IN7(na21_2),
                      .IN8(na58_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x30y77     80'h00_0018_00_0040_0AF7_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1028_1 ( .OUT(na1028_1), .IN1(1'b1), .IN2(~na871_2), .IN3(1'b1), .IN4(na1703_2), .IN5(~na611_1), .IN6(~na20_2), .IN7(~na21_2),
                      .IN8(na1702_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///ICOMP/      x32y75     80'h00_0060_00_0000_0C08_FFC9
C_ICOMP    #(.CPE_CFG (9'b0_1000_0000)) 
           _a1029_4 ( .OUT(na1029_2), .IN1(na1745_2), .IN2(na613_1), .IN3(1'b1), .IN4(na22_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x32y76     80'h00_0018_00_0040_0A99_0033
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1030_1 ( .OUT(na1030_1), .IN1(1'b1), .IN2(~na871_2), .IN3(1'b1), .IN4(~na1703_2), .IN5(~na57_1), .IN6(1'b0), .IN7(1'b0),
                      .IN8(~na58_2), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1031 ( .O(ant_433mhz), .A(na1602_10) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000010)) 
           _a1032 ( .Y(na1032_1), .I(btn) );
CPE_IBF    #(.BUF_CFG (72'h000001000000000090)) 
           _a1033 ( .Y(na1033_1), .I(clk_10mhz) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1034 ( .O(led), .A(na1603_10) );
CPE_OBF    #(.BUF_CFG (72'h000000000100010900)) 
           _a1035 ( .O(wifi_gpio0), .A(na1604_10) );
// C_/C_0_1///      x47y55     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1036_2 ( .OUT(na1036_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1036_6 ( .COUTY1(na1036_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1036_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_/C_0_1///      x54y69     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1037_2 ( .OUT(na1037_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1037_6 ( .COUTY1(na1037_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1037_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_05_08_0A_20_82)) 
           _a1038 ( .USR_PLL_LOCKED_STDY(_d6), .USR_PLL_LOCKED(_d7), .CLK270(na1038_3), .CLK180(na1038_4), .CLK90(na1038_5), .CLK0(na1038_6),
                    .CLK_REF_OUT(_d8), .CLK_REF(na1040_1), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
CC_PLL     #(.PLL_CFG (96'h01_CB_01_10_64_00_04_01_08_08_30_82)) 
           _a1039 ( .USR_PLL_LOCKED_STDY(_d9), .USR_PLL_LOCKED(_d10), .CLK270(na1039_3), .CLK180(na1039_4), .CLK90(na1039_5), .CLK0(na1039_6),
                    .CLK_REF_OUT(_d11), .CLK_REF(na1040_2), .CLK_FEEDBACK(1'b0), .USR_CLK_REF(1'b0), .USR_LOCKED_STDY_RST(1'b0), .USR_SET_SEL(1'b0) );
CLKIN      #(.CLKIN_CFG (32'h0000_0000)) 
           _a1040 ( .PCLK0(na1040_1), .PCLK1(na1040_2), .PCLK2(_d12), .PCLK3(_d13), .CLK0(na1033_1), .CLK1(1'b0), .CLK2(1'b0), .CLK3(1'b0),
                    .SER_CLK(1'b0), .SPI_CLK(1'b0), .JTAG_CLK(1'b0) );
// C_///AND/      x27y75     80'h00_0060_00_0000_0C08_FF3C
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1041_4 ( .OUT(na1041_2), .IN1(1'b1), .IN2(na98_2), .IN3(1'b1), .IN4(~na99_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x27y76     80'h00_0018_00_0000_0C66_CC00
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1042_1 ( .OUT(na1042_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na98_2), .IN7(1'b0), .IN8(na99_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x19y73     80'h00_0060_00_0000_0C08_FFAC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1043_4 ( .OUT(na1043_2), .IN1(1'b1), .IN2(na98_2), .IN3(na1640_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x22y74     80'h00_0018_00_0000_0C88_53FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1044_1 ( .OUT(na1044_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na98_2), .IN7(~na1640_2), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x30y75     80'h00_0060_00_0000_0C08_FFC3
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1045_4 ( .OUT(na1045_2), .IN1(1'b1), .IN2(~na98_1), .IN3(1'b1), .IN4(na99_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x19y77     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1046_1 ( .OUT(na1046_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1643_2), .IN6(1'b1), .IN7(1'b1), .IN8(~na99_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x22y78     80'h00_0060_00_0000_0C08_FFC5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1047_4 ( .OUT(na1047_2), .IN1(~na1643_2), .IN2(1'b1), .IN3(1'b1), .IN4(na99_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x26y80     80'h00_0018_00_0000_0C88_33FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1048_1 ( .OUT(na1048_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na98_1), .IN7(1'b1), .IN8(~na99_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x22y73     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1049_4 ( .OUT(na1049_2), .IN1(1'b1), .IN2(na98_1), .IN3(1'b1), .IN4(na99_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_/C_0_1///      x53y67     80'h00_CF00_12_0800_0C00_FFFF
C_C_0_1    #(.CPE_CFG (9'bX_0000_0000)) 
           _a1050_2 ( .OUT(na1050_1), .CLK(1'b1), .EN(1'b1), .SR(1'b0), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN() );
C_CPlines  #(.CPE_CFG (19'h1_2080)) 
           _a1050_6 ( .COUTY1(na1050_4), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(na1050_1),
                      .OUT2(1'b0), .COMP_OUT(1'b0) );
// C_Route1////      x35y77     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a1051_1 ( .OUT(na1051_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na580_4), .PINX(1'b0), .PINY1(1'b0) );
// C_Route1////      x26y76     80'h00_0018_00_0050_0C66_0000
C_Route1   #(.CPE_CFG (9'b0_0001_0000)) 
           _a1052_1 ( .OUT(na1052_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na620_4), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x29y76     80'h00_0018_00_0000_0C88_C3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1054_1 ( .OUT(na1054_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na98_2), .IN7(1'b1), .IN8(na99_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x27y79     80'h00_0060_00_0000_0C06_FFCC
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1055_4 ( .OUT(na1055_2), .IN1(1'b0), .IN2(na98_1), .IN3(1'b0), .IN4(na99_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4a////      x29y81     80'h00_0018_00_0040_0CE8_C300
C_MX4a     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1056_1 ( .OUT(na1056_1), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(~na99_2), .IN5(1'b1), .IN6(~na98_2), .IN7(1'b1), .IN8(na99_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x58y70     80'h00_0018_00_0040_0A61_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1060_1 ( .OUT(na1060_1), .IN1(1'b1), .IN2(na1776_2), .IN3(1'b1), .IN4(na116_2), .IN5(1'b1), .IN6(na1779_2), .IN7(na969_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y75     80'h00_0018_00_0040_0A92_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1061_1 ( .OUT(na1061_1), .IN1(1'b1), .IN2(~na891_1), .IN3(na1649_2), .IN4(1'b1), .IN5(na895_1), .IN6(1'b1), .IN7(1'b0), .IN8(na1750_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x61y75     80'h00_0018_00_0040_0A92_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1062_1 ( .OUT(na1062_1), .IN1(1'b1), .IN2(~na1778_2), .IN3(na111_1), .IN4(1'b1), .IN5(na1780_2), .IN6(1'b1), .IN7(1'b0),
                      .IN8(na971_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x49y68     80'h00_0018_00_0040_0A92_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1063_1 ( .OUT(na1063_1), .IN1(1'b1), .IN2(~na893_1), .IN3(na112_1), .IN4(1'b1), .IN5(na897_1), .IN6(1'b1), .IN7(1'b0), .IN8(na1752_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y73     80'h00_0018_00_0040_0A61_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1064_1 ( .OUT(na1064_1), .IN1(1'b1), .IN2(na1779_2), .IN3(1'b1), .IN4(na113_2), .IN5(1'b1), .IN6(na1770_2), .IN7(na958_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y77     80'h00_0018_00_0040_0A61_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1065_1 ( .OUT(na1065_1), .IN1(na1646_2), .IN2(1'b1), .IN3(1'b1), .IN4(na1750_2), .IN5(1'b1), .IN6(na899_1), .IN7(na1754_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y79     80'h00_0018_00_0040_0A92_00A3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1066_1 ( .OUT(na1066_1), .IN1(1'b1), .IN2(~na1781_2), .IN3(na115_2), .IN4(1'b1), .IN5(na1771_2), .IN6(1'b1), .IN7(1'b0),
                      .IN8(na960_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x60y71     80'h00_0018_00_0040_0A92_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1067_1 ( .OUT(na1067_1), .IN1(~na981_1), .IN2(1'b1), .IN3(1'b1), .IN4(na116_2), .IN5(na985_1), .IN6(1'b1), .IN7(1'b0), .IN8(na1795_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x53y65     80'h00_0018_00_0040_0A61_00CA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1068_1 ( .OUT(na1068_1), .IN1(na118_1), .IN2(1'b1), .IN3(1'b1), .IN4(na723_2), .IN5(1'b1), .IN6(na727_2), .IN7(na1711_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x57y71     80'h00_0018_00_0040_0A61_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1069_1 ( .OUT(na1069_1), .IN1(1'b1), .IN2(na983_1), .IN3(na111_1), .IN4(1'b1), .IN5(1'b1), .IN6(na987_1), .IN7(na1797_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y66     80'h00_0018_00_0040_0A61_00AA
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1070_1 ( .OUT(na1070_1), .IN1(na1708_2), .IN2(1'b1), .IN3(na112_1), .IN4(1'b1), .IN5(1'b1), .IN6(na729_2), .IN7(na1713_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x55y75     80'h00_0018_00_0040_0A92_00C5
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1071_1 ( .OUT(na1071_1), .IN1(~na985_1), .IN2(1'b1), .IN3(1'b1), .IN4(na113_2), .IN5(na974_1), .IN6(1'b1), .IN7(1'b0), .IN8(na1784_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x50y70     80'h00_0018_00_0040_0A61_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1072_1 ( .OUT(na1072_1), .IN1(1'b1), .IN2(na727_2), .IN3(1'b1), .IN4(na114_1), .IN5(1'b1), .IN6(na1717_2), .IN7(na731_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x59y67     80'h00_0018_00_0040_0A61_00AC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1073_1 ( .OUT(na1073_1), .IN1(1'b1), .IN2(na987_1), .IN3(na115_2), .IN4(1'b1), .IN5(1'b1), .IN6(na976_1), .IN7(na1786_2),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x49y63     80'h00_0018_00_0000_0C88_F4FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1075_1 ( .OUT(na1075_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1578_1), .IN6(na844_2), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x50y66     80'h00_0060_00_0000_0C06_FF09
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1076_4 ( .OUT(na1076_2), .IN1(na1578_1), .IN2(~na844_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x53y60     80'h00_0018_00_0040_0A32_000C
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1079_1 ( .OUT(na1079_1), .IN1(1'b1), .IN2(na1652_2), .IN3(1'b0), .IN4(1'b0), .IN5(na165_1), .IN6(~na553_1), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y59     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1080_1 ( .OUT(na1080_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na182_1), .IN5(1'b0), .IN6(~na553_2), .IN7(1'b0), .IN8(~na1016_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x50y60     80'h00_0018_00_0040_0A33_0003
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1081_1 ( .OUT(na1081_1), .IN1(1'b1), .IN2(~na1652_2), .IN3(1'b0), .IN4(1'b0), .IN5(~na555_1), .IN6(~na1019_1), .IN7(1'b0),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x48y57     80'h00_0018_00_0040_0A55_0030
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1082_1 ( .OUT(na1082_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b1), .IN4(~na182_1), .IN5(~na555_2), .IN6(1'b0), .IN7(~na1022_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x53y59     80'h00_0018_00_0040_0AAA_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1083_1 ( .OUT(na1083_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na182_1), .IN5(1'b0), .IN6(~na557_1), .IN7(1'b0), .IN8(~na1024_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX2b////      x43y50     80'h00_0018_00_0040_0AA2_003F
C_MX2b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1084_1 ( .OUT(na1084_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(~na182_1), .IN5(1'b0), .IN6(~na557_2), .IN7(1'b0), .IN8(na90_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x39y74     80'h00_0018_00_0040_0A61_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1085_1 ( .OUT(na1085_1), .IN1(1'b1), .IN2(na234_2), .IN3(1'b1), .IN4(na235_1), .IN5(1'b1), .IN6(na1634_2), .IN7(na46_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x37y70     80'h00_0018_00_0000_0C88_5AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1087_1 ( .OUT(na1087_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na47_1), .IN6(1'b1), .IN7(~na46_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x40y74     80'h00_0018_00_0040_0A92_00C3
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1088_1 ( .OUT(na1088_1), .IN1(1'b1), .IN2(~na234_2), .IN3(1'b1), .IN4(na235_1), .IN5(na47_1), .IN6(1'b1), .IN7(1'b0), .IN8(na1635_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x35y73     80'h00_0060_00_0000_0C08_FFA5
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1090_4 ( .OUT(na1090_2), .IN1(~na47_1), .IN2(1'b1), .IN3(na48_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_MX4b////      x40y76     80'h00_0018_00_0040_0A61_00CC
C_MX4b     #(.CPE_CFG (9'b0_0000_0000)) 
           _a1091_1 ( .OUT(na1091_1), .IN1(1'b1), .IN2(na234_2), .IN3(1'b1), .IN4(na235_1), .IN5(1'b1), .IN6(na1636_2), .IN7(na48_1),
                      .IN8(1'b0), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x50y68     80'h00_0078_00_0000_0C66_C99A
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1092_1 ( .OUT(na1092_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na722_2), .IN6(~na269_1), .IN7(1'b0), .IN8(na176_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1092_4 ( .OUT(na1092_2), .IN1(na1075_1), .IN2(1'b0), .IN3(na721_1), .IN4(~na176_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x55y63     80'h00_0078_00_0000_0C66_A965
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1095_1 ( .OUT(na1095_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na724_1), .IN6(~na279_1), .IN7(na275_2), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1095_4 ( .OUT(na1095_2), .IN1(~na274_1), .IN2(1'b0), .IN3(na275_1), .IN4(na723_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR////      x34y70     80'h00_0018_00_0000_0666_95C3
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1097_1 ( .OUT(na1097_1), .IN1(1'b0), .IN2(~na1025_1), .IN3(1'b0), .IN4(na184_1), .IN5(~na40_1), .IN6(1'b0), .IN7(na185_2),
                      .IN8(~na181_1), .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x59y75     80'h00_0078_00_0000_0C66_AA56
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1098_1 ( .OUT(na1098_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1769_2), .IN6(1'b0), .IN7(na962_1), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1098_4 ( .OUT(na1098_2), .IN1(na1769_2), .IN2(na295_1), .IN3(~na962_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x55y81     80'h00_0018_00_0000_0C88_A3FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1100_1 ( .OUT(na1100_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(~na1770_2), .IN7(na962_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x58y68     80'h00_0060_00_0000_0C06_FF9C
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1102_4 ( .OUT(na1102_2), .IN1(1'b0), .IN2(na1779_2), .IN3(na965_1), .IN4(~na116_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x58y81     80'h00_0078_00_0000_0C88_CCCC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1112_1 ( .OUT(na1112_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na1775_2), .IN7(1'b1), .IN8(na960_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1112_4 ( .OUT(na1112_2), .IN1(1'b1), .IN2(na899_1), .IN3(1'b1), .IN4(na963_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND/      x56y80     80'h00_0060_00_0000_0C08_FFCC
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1113_4 ( .OUT(na1113_2), .IN1(1'b1), .IN2(na901_1), .IN3(1'b1), .IN4(na963_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_XOR///XOR/      x55y77     80'h00_0078_00_0000_0C66_0665
C_XOR      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1114_1 ( .OUT(na1114_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na978_1), .IN6(na1782_2), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1114_4 ( .OUT(na1114_2), .IN1(~na978_1), .IN2(1'b0), .IN3(na1783_2), .IN4(na321_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x60y80     80'h00_0018_00_0000_0C88_3AFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1116_1 ( .OUT(na1116_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na978_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1784_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///XOR/      x55y70     80'h00_0060_00_0000_0C06_FF9A
C_XOR      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1118_4 ( .OUT(na1118_2), .IN1(na981_1), .IN2(1'b0), .IN3(na1794_2), .IN4(~na116_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND///AND/      x57y77     80'h00_0078_00_0000_0C88_CCAC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1128_1 ( .OUT(na1128_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na976_1), .IN7(1'b1), .IN8(na1789_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1128_4 ( .OUT(na1128_2), .IN1(1'b1), .IN2(na979_1), .IN3(na731_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND////      x55y78     80'h00_0018_00_0000_0C88_CCFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1129_1 ( .OUT(na1129_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na979_1), .IN7(1'b1), .IN8(na733_2),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_///AND*/      x26y40     80'h00_0060_00_0000_0C07_FFF0
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1130_4 ( .OUT(na1130_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND//O_0/AND/      x26y41     80'h00_0078_09_6000_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1131_1 ( .OUT(na1131_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a1131_3 ( .COMP_OUT(na1131_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1131_4 ( .OUT(na1131_2), .IN1(1'b1), .IN2(na663_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1131_6 ( .COUTX(na1131_3), .POUTX(na1131_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1131_1), .OUT2(na1131_2), .COMP_OUT(na1131_3_i) );
// C_AND*/D//AND*/D      x26y42     80'h00_FE00_89_6000_0387_FAFC
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1132_1 ( .OUT(na1132_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na251_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1132_2 ( .OUT(na1132_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1132_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1132_4 ( .OUT(na1132_2_i), .IN1(1'b1), .IN2(na634_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1132_5 ( .OUT(na1132_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1132_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1132_6 ( .COUTX(na1132_3), .POUTX(na1132_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1132_1), .OUT2(na1132_2), .COMP_OUT(1'b0) );
// C_AND/D//AND/D      x26y43     80'h00_FE00_89_6000_0C88_FCAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1133_1 ( .OUT(na1133_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na635_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1133_2 ( .OUT(na1133_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1133_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1133_4 ( .OUT(na1133_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na636_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1133_5 ( .OUT(na1133_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1133_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1133_6 ( .COUTX(na1133_3), .POUTX(na1133_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1133_1), .OUT2(na1133_2), .COMP_OUT(1'b0) );
// C_AND*/D//AND*/D      x26y44     80'h00_FE00_89_6000_0387_CFCF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1134_1 ( .OUT(na1134_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na480_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1134_2 ( .OUT(na1134_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1134_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1134_4 ( .OUT(na1134_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na638_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1134_5 ( .OUT(na1134_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1134_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1134_6 ( .COUTX(na1134_3), .POUTX(na1134_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1134_1), .OUT2(na1134_2), .COMP_OUT(1'b0) );
// C_AND/D//AND/D      x26y45     80'h00_FE00_89_6000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1135_1 ( .OUT(na1135_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na489_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1135_2 ( .OUT(na1135_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1135_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1135_4 ( .OUT(na1135_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na640_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1135_5 ( .OUT(na1135_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1135_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1135_6 ( .COUTX(na1135_3), .POUTX(na1135_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1135_1), .OUT2(na1135_2), .COMP_OUT(1'b0) );
// C_AND*/D//AND*/D      x26y46     80'h00_FE00_89_6000_0387_CFAF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1136_1 ( .OUT(na1136_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na491_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1136_2 ( .OUT(na1136_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1136_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1136_4 ( .OUT(na1136_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na642_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1136_5 ( .OUT(na1136_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1136_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1136_6 ( .COUTX(na1136_3), .POUTX(na1136_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1136_1), .OUT2(na1136_2), .COMP_OUT(1'b0) );
// C_AND/D//AND/D      x26y47     80'h00_FE00_89_6000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1137_1 ( .OUT(na1137_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na493_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1137_2 ( .OUT(na1137_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1137_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1137_4 ( .OUT(na1137_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na644_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1137_5 ( .OUT(na1137_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1137_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1137_6 ( .COUTX(na1137_3), .POUTX(na1137_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1137_1), .OUT2(na1137_2), .COMP_OUT(1'b0) );
// C_AND*/D//AND*/D      x26y48     80'h00_FE00_89_6000_0387_CFAF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1138_1 ( .OUT(na1138_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na495_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1138_2 ( .OUT(na1138_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1138_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1138_4 ( .OUT(na1138_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na646_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1138_5 ( .OUT(na1138_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1138_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1138_6 ( .COUTX(na1138_3), .POUTX(na1138_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1138_1), .OUT2(na1138_2), .COMP_OUT(1'b0) );
// C_AND/D//AND/D      x26y49     80'h00_FE00_89_6000_0C88_AFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1139_1 ( .OUT(na1139_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na471_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1139_2 ( .OUT(na1139_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1139_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1139_4 ( .OUT(na1139_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na648_2), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1139_5 ( .OUT(na1139_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1139_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1139_6 ( .COUTX(na1139_3), .POUTX(na1139_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1139_1), .OUT2(na1139_2), .COMP_OUT(1'b0) );
// C_AND*/D//AND*/D      x26y50     80'h00_FE00_89_6000_0387_CFCF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1140_1 ( .OUT(na1140_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na473_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1140_2 ( .OUT(na1140_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1140_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1140_4 ( .OUT(na1140_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na650_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1140_5 ( .OUT(na1140_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1140_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1140_6 ( .COUTX(na1140_3), .POUTX(na1140_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1140_1), .OUT2(na1140_2), .COMP_OUT(1'b0) );
// C_AND/D//AND/D      x26y51     80'h00_FE00_89_6000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1141_1 ( .OUT(na1141_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na475_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1141_2 ( .OUT(na1141_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1141_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1141_4 ( .OUT(na1141_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na652_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1141_5 ( .OUT(na1141_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1141_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1141_6 ( .COUTX(na1141_3), .POUTX(na1141_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1141_1), .OUT2(na1141_2), .COMP_OUT(1'b0) );
// C_AND*/D//AND*/D      x26y52     80'h00_FE00_89_6000_0387_CFAF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1142_1 ( .OUT(na1142_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na477_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1142_2 ( .OUT(na1142_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1142_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1142_4 ( .OUT(na1142_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na654_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1142_5 ( .OUT(na1142_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1142_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1142_6 ( .COUTX(na1142_3), .POUTX(na1142_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1142_1), .OUT2(na1142_2), .COMP_OUT(1'b0) );
// C_AND/D//AND/D      x26y53     80'h00_FE00_89_6000_0C88_AFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1143_1 ( .OUT(na1143_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na479_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1143_2 ( .OUT(na1143_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1143_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1143_4 ( .OUT(na1143_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(na656_2), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1143_5 ( .OUT(na1143_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1143_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1143_6 ( .COUTX(na1143_3), .POUTX(na1143_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1143_1), .OUT2(na1143_2), .COMP_OUT(1'b0) );
// C_AND*/D//AND*/D      x26y54     80'h00_FE00_89_6000_0387_CFFA
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1144_1 ( .OUT(na1144_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na482_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1144_2 ( .OUT(na1144_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1144_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1144_4 ( .OUT(na1144_2_i), .IN1(na658_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1144_5 ( .OUT(na1144_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1144_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1144_6 ( .COUTX(na1144_3), .POUTX(na1144_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1144_1), .OUT2(na1144_2), .COMP_OUT(1'b0) );
// C_AND/D//AND/D      x26y55     80'h00_FE00_89_6000_0C88_AFFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1145_1 ( .OUT(na1145_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(na484_1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1145_2 ( .OUT(na1145_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1145_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1145_4 ( .OUT(na1145_2_i), .IN1(na660_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1145_5 ( .OUT(na1145_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1145_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1145_6 ( .COUTX(na1145_3), .POUTX(na1145_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1145_1), .OUT2(na1145_2), .COMP_OUT(1'b0) );
// C_AND*/D//AND*/D      x26y56     80'h00_FE00_89_6000_0387_CFCF
C_AND      #(.CPE_CFG (9'b1_0000_0000)) 
           _a1146_1 ( .OUT(na1146_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na486_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1146_2 ( .OUT(na1146_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1146_1_i) );
C_AND      #(.CPE_CFG (9'b1_1000_0000)) 
           _a1146_4 ( .OUT(na1146_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na662_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1146_5 ( .OUT(na1146_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1146_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1146_6 ( .COUTX(na1146_3), .POUTX(na1146_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1146_1), .OUT2(na1146_2), .COMP_OUT(1'b0) );
// C_AND/D//AND/D      x26y57     80'h00_FE00_89_6000_0C88_CFCF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1147_1 ( .OUT(na1147_1_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na662_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0000)) 
           _a1147_2 ( .OUT(na1147_1), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1147_1_i) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1147_4 ( .OUT(na1147_2_i), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(na662_1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_D        #(.CPE_CFG (9'bX_0000_0100)) 
           _a1147_5 ( .OUT(na1147_2), .CLK(na624_2), .EN(1'b1), .SR(1'b1), .CINY2(1'b0), .PINY2(1'b0), .RAM_I(1'b0), .CP_O(1'b0), .D_IN(na1147_2_i) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1147_6 ( .COUTX(na1147_3), .POUTX(na1147_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1147_1), .OUT2(na1147_2), .COMP_OUT(1'b0) );
// C_AND///AND/      x27y37     80'h00_0078_12_0000_0C88_FFF0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1148_1 ( .OUT(na1148_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1148_4 ( .OUT(na1148_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1148_6 ( .COUTY1(na1148_4), .POUTY1(na1148_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1148_1), .OUT2(na1148_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x27y38     80'h00_0018_04_2056_5888_0CC0
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1149_1 ( .OUT(na1149_1), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1148_4), .PINX(1'b0), .PINY1(na1148_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1149_3 ( .COMP_OUT(na1149_3_i), .COMB1(na1149_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1149_6 ( .COUTY1(na1149_4), .COUTY2(na1149_5), .POUTY1(na1149_7), .CINX(1'b0), .CINY1(na1148_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1148_7), .PINY2(1'b0), .OUT1(na1149_1), .OUT2(1'b0), .COMP_OUT(na1149_3_i) );
// C_MULTFa//O_O2//      x27y39     80'h00_0018_13_A477_34A6_0C0C
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1150_1 ( .COUTX(na1150_3), .COUTY1(na1150_4), .COUTY2(na1150_5), .POUTY1(na1150_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1149_4),
                      .CINY2(na1149_5), .PINX(1'b0), .PINY1(na1149_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x27y40     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1151_1 ( .OUT(na1151_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1150_4), .PINX(1'b0), .PINY1(na1150_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1151_3 ( .COMP_OUT(na1151_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1151_4 ( .OUT(na1151_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1150_4), .PINX(1'b0), .PINY1(na1150_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1151_6 ( .COUTX(na1151_3), .COUTY1(na1151_4), .COUTY2(na1151_5), .POUTY1(na1151_7), .POUTY2(na1151_8), .CINX(1'b0), .CINY1(na1150_4),
                      .CINY2(na1150_5), .PINX(1'b0), .PINY1(na1150_7), .PINY2(1'b0), .OUT1(na1151_1), .OUT2(na1151_2), .COMP_OUT(na1151_3_i) );
// C_MULT///MULT/      x27y41     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1152_1 ( .COUTY1(na1152_4), .COUTY2(na1152_5), .POUTY1(na1152_7), .POUTY2(na1152_8), .IN1(na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(1'b0),
                      .CINY1(na1151_4), .CINY2(na1151_5), .PINX(1'b0), .PINY1(na1151_7), .PINY2(na1151_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y42     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1153_1 ( .COUTX(na1153_3), .COUTY1(na1153_4), .COUTY2(na1153_5), .POUTX(na1153_6), .POUTY1(na1153_7), .POUTY2(na1153_8),
                      .IN1(~na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1152_4), .CINY2(na1152_5), .PINX(1'b0), .PINY1(na1152_7), .PINY2(na1152_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y43     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1154_1 ( .COUTX(na1154_3), .COUTY1(na1154_4), .COUTY2(na1154_5), .POUTX(na1154_6), .POUTY1(na1154_7), .POUTY2(na1154_8),
                      .IN1(na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1153_4), .CINY2(na1153_5), .PINX(1'b0), .PINY1(na1153_7), .PINY2(na1153_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y44     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1155_1 ( .COUTX(na1155_3), .COUTY1(na1155_4), .COUTY2(na1155_5), .POUTX(na1155_6), .POUTY1(na1155_7), .POUTY2(na1155_8),
                      .IN1(~na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1154_4), .CINY2(na1154_5), .PINX(1'b0), .PINY1(na1154_7), .PINY2(na1154_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y45     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1156_1 ( .COUTX(na1156_3), .COUTY1(na1156_4), .COUTY2(na1156_5), .POUTX(na1156_6), .POUTY1(na1156_7), .POUTY2(na1156_8),
                      .IN1(na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1155_4), .CINY2(na1155_5), .PINX(1'b0), .PINY1(na1155_7), .PINY2(na1155_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y46     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1157_1 ( .COUTX(na1157_3), .COUTY1(na1157_4), .COUTY2(na1157_5), .POUTX(na1157_6), .POUTY1(na1157_7), .POUTY2(na1157_8),
                      .IN1(~na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1156_4), .CINY2(na1156_5), .PINX(1'b0), .PINY1(na1156_7), .PINY2(na1156_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y47     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1158_1 ( .COUTX(na1158_3), .COUTY1(na1158_4), .COUTY2(na1158_5), .POUTX(na1158_6), .POUTY1(na1158_7), .POUTY2(na1158_8),
                      .IN1(na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1157_4), .CINY2(na1157_5), .PINX(1'b0), .PINY1(na1157_7), .PINY2(na1157_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y48     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1159_1 ( .COUTX(na1159_3), .COUTY1(na1159_4), .COUTY2(na1159_5), .POUTX(na1159_6), .POUTY1(na1159_7), .POUTY2(na1159_8),
                      .IN1(~na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1158_4), .CINY2(na1158_5), .PINX(1'b0), .PINY1(na1158_7), .PINY2(na1158_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y49     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1160_1 ( .COUTX(na1160_3), .COUTY1(na1160_4), .COUTY2(na1160_5), .POUTX(na1160_6), .POUTY1(na1160_7), .POUTY2(na1160_8),
                      .IN1(na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1159_4), .CINY2(na1159_5), .PINX(1'b0), .PINY1(na1159_7), .PINY2(na1159_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y50     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1161_1 ( .COUTX(na1161_3), .COUTY1(na1161_4), .COUTY2(na1161_5), .POUTX(na1161_6), .POUTY1(na1161_7), .POUTY2(na1161_8),
                      .IN1(~na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1160_4), .CINY2(na1160_5), .PINX(1'b0), .PINY1(na1160_7), .PINY2(na1160_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y51     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1162_1 ( .COUTX(na1162_3), .COUTY1(na1162_4), .COUTY2(na1162_5), .POUTX(na1162_6), .POUTY1(na1162_7), .POUTY2(na1162_8),
                      .IN1(na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1161_4), .CINY2(na1161_5), .PINX(1'b0), .PINY1(na1161_7), .PINY2(na1161_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y52     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1163_1 ( .COUTX(na1163_3), .COUTY1(na1163_4), .COUTY2(na1163_5), .POUTX(na1163_6), .POUTY1(na1163_7), .POUTY2(na1163_8),
                      .IN1(~na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1162_4), .CINY2(na1162_5), .PINX(1'b0), .PINY1(na1162_7), .PINY2(na1162_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1164_1 ( .COUTX(na1164_3), .COUTY1(na1164_4), .COUTY2(na1164_5), .POUTX(na1164_6), .POUTY1(na1164_7), .POUTY2(na1164_8),
                      .IN1(na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1163_4), .CINY2(na1163_5), .PINX(1'b0), .PINY1(na1163_7), .PINY2(na1163_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1165_1 ( .COUTX(na1165_3), .COUTY1(na1165_4), .COUTY2(na1165_5), .POUTX(na1165_6), .POUTY1(na1165_7), .POUTY2(na1165_8),
                      .IN1(~na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1164_4), .CINY2(na1164_5), .PINX(1'b0), .PINY1(na1164_7), .PINY2(na1164_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1166_1 ( .COUTX(na1166_3), .COUTY1(na1166_4), .COUTY2(na1166_5), .POUTX(na1166_6), .POUTY1(na1166_7), .POUTY2(na1166_8),
                      .IN1(na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1165_4), .CINY2(na1165_5), .PINX(1'b0), .PINY1(na1165_7), .PINY2(na1165_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1167_1 ( .COUTX(na1167_3), .COUTY1(na1167_4), .COUTY2(na1167_5), .POUTX(na1167_6), .POUTY1(na1167_7), .POUTY2(na1167_8),
                      .IN1(~na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1166_4), .CINY2(na1166_5), .PINX(1'b0), .PINY1(na1166_7), .PINY2(na1166_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x27y57     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1168_1 ( .COUTX(na1168_3), .COUTY1(na1168_4), .COUTY2(na1168_5), .POUTX(na1168_6), .POUTY1(na1168_7), .POUTY2(na1168_8),
                      .IN1(na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1167_4), .CINY2(na1167_5), .PINX(1'b0), .PINY1(na1167_7), .PINY2(na1167_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x27y58     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1169_3 ( .COMP_OUT(na1169_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1169_4 ( .OUT(na1169_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1168_4), .PINX(1'b0), .PINY1(na1168_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1169_6 ( .COUTX(na1169_3), .POUTX(na1169_6), .CINX(1'b0), .CINY1(na1168_4), .CINY2(na1168_5), .PINX(1'b0), .PINY1(na1168_7),
                      .PINY2(na1168_8), .OUT1(1'b0), .OUT2(na1169_2), .COMP_OUT(na1169_3_i) );
// C_AND///AND/      x28y38     80'h00_0078_12_0000_0C88_FFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1170_1 ( .OUT(na1170_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1170_4 ( .OUT(na1170_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1170_6 ( .COUTY1(na1170_4), .POUTY1(na1170_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1170_1), .OUT2(na1170_2), .COMP_OUT(1'b0) );
// C_OR//O_O1//      x28y39     80'h00_0018_04_2056_5EEE_0CC0
C_OR       #(.CPE_CFG (9'b0_0001_0110)) 
           _a1171_1 ( .OUT(na1171_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(na1150_3), .CINY1(na1170_4), .PINX(1'b0), .PINY1(na1170_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1171_3 ( .COMP_OUT(na1171_3_i), .COMB1(na1171_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1171_6 ( .COUTY1(na1171_4), .COUTY2(na1171_5), .POUTY1(na1171_7), .CINX(na1150_3), .CINY1(na1170_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1170_7), .PINY2(1'b0), .OUT1(na1171_1), .OUT2(1'b0), .COMP_OUT(na1171_3_i) );
// C_MULTFb//O_O2//      x28y40     80'h00_0018_13_A477_3EA6_0CCC
C_MULTFb   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1172_1 ( .COUTX(na1172_3), .COUTY1(na1172_4), .COUTY2(na1172_5), .POUTY1(na1172_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1151_3), .CINY1(na1171_4),
                      .CINY2(na1171_5), .PINX(1'b0), .PINY1(na1171_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_O2/AND/      x28y41     80'h00_0078_35_A471_3C88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1173_1 ( .OUT(na1173_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1172_4), .PINX(1'b0), .PINY1(na1172_7) );
C_O_O2     #(.CPE_CFG ()) 
           _a1173_3 ( .COMP_OUT(na1173_3_i), .COMB1(1'b0), .COMB2(na1173_2) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1173_4 ( .OUT(na1173_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1172_4), .PINX(1'b0), .PINY1(na1172_7) );
C_CPlines  #(.CPE_CFG (19'h3_5A47)) 
           _a1173_6 ( .COUTX(na1173_3), .COUTY1(na1173_4), .COUTY2(na1173_5), .POUTY1(na1173_7), .POUTY2(na1173_8), .CINX(1'b0), .CINY1(na1172_4),
                      .CINY2(na1172_5), .PINX(1'b0), .PINY1(na1172_7), .PINY2(1'b0), .OUT1(na1173_1), .OUT2(na1173_2), .COMP_OUT(na1173_3_i) );
// C_MULT///MULT/      x28y42     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1174_1 ( .COUTY1(na1174_4), .COUTY2(na1174_5), .POUTY1(na1174_7), .POUTY2(na1174_8), .IN1(~na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1153_3),
                      .CINY1(na1173_4), .CINY2(na1173_5), .PINX(na1153_6), .PINY1(na1173_7), .PINY2(na1173_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y43     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1175_1 ( .COUTX(na1175_3), .COUTY1(na1175_4), .COUTY2(na1175_5), .POUTX(na1175_6), .POUTY1(na1175_7), .POUTY2(na1175_8),
                      .IN1(na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1154_3), .CINY1(na1174_4), .CINY2(na1174_5), .PINX(na1154_6), .PINY1(na1174_7), .PINY2(na1174_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y44     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1176_1 ( .COUTX(na1176_3), .COUTY1(na1176_4), .COUTY2(na1176_5), .POUTX(na1176_6), .POUTY1(na1176_7), .POUTY2(na1176_8),
                      .IN1(~na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1155_3), .CINY1(na1175_4), .CINY2(na1175_5), .PINX(na1155_6), .PINY1(na1175_7), .PINY2(na1175_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y45     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1177_1 ( .COUTX(na1177_3), .COUTY1(na1177_4), .COUTY2(na1177_5), .POUTX(na1177_6), .POUTY1(na1177_7), .POUTY2(na1177_8),
                      .IN1(na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1156_3), .CINY1(na1176_4), .CINY2(na1176_5), .PINX(na1156_6), .PINY1(na1176_7), .PINY2(na1176_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y46     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1178_1 ( .COUTX(na1178_3), .COUTY1(na1178_4), .COUTY2(na1178_5), .POUTX(na1178_6), .POUTY1(na1178_7), .POUTY2(na1178_8),
                      .IN1(~na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1157_3), .CINY1(na1177_4), .CINY2(na1177_5), .PINX(na1157_6), .PINY1(na1177_7), .PINY2(na1177_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y47     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1179_1 ( .COUTX(na1179_3), .COUTY1(na1179_4), .COUTY2(na1179_5), .POUTX(na1179_6), .POUTY1(na1179_7), .POUTY2(na1179_8),
                      .IN1(na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1158_3), .CINY1(na1178_4), .CINY2(na1178_5), .PINX(na1158_6), .PINY1(na1178_7), .PINY2(na1178_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y48     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1180_1 ( .COUTX(na1180_3), .COUTY1(na1180_4), .COUTY2(na1180_5), .POUTX(na1180_6), .POUTY1(na1180_7), .POUTY2(na1180_8),
                      .IN1(~na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1159_3), .CINY1(na1179_4), .CINY2(na1179_5), .PINX(na1159_6), .PINY1(na1179_7), .PINY2(na1179_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y49     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1181_1 ( .COUTX(na1181_3), .COUTY1(na1181_4), .COUTY2(na1181_5), .POUTX(na1181_6), .POUTY1(na1181_7), .POUTY2(na1181_8),
                      .IN1(na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1160_3), .CINY1(na1180_4), .CINY2(na1180_5), .PINX(na1160_6), .PINY1(na1180_7), .PINY2(na1180_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y50     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1182_1 ( .COUTX(na1182_3), .COUTY1(na1182_4), .COUTY2(na1182_5), .POUTX(na1182_6), .POUTY1(na1182_7), .POUTY2(na1182_8),
                      .IN1(~na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1161_3), .CINY1(na1181_4), .CINY2(na1181_5), .PINX(na1161_6), .PINY1(na1181_7), .PINY2(na1181_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y51     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1183_1 ( .COUTX(na1183_3), .COUTY1(na1183_4), .COUTY2(na1183_5), .POUTX(na1183_6), .POUTY1(na1183_7), .POUTY2(na1183_8),
                      .IN1(na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1162_3), .CINY1(na1182_4), .CINY2(na1182_5), .PINX(na1162_6), .PINY1(na1182_7), .PINY2(na1182_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y52     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1184_1 ( .COUTX(na1184_3), .COUTY1(na1184_4), .COUTY2(na1184_5), .POUTX(na1184_6), .POUTY1(na1184_7), .POUTY2(na1184_8),
                      .IN1(~na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1163_3), .CINY1(na1183_4), .CINY2(na1183_5), .PINX(na1163_6), .PINY1(na1183_7), .PINY2(na1183_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1185_1 ( .COUTX(na1185_3), .COUTY1(na1185_4), .COUTY2(na1185_5), .POUTX(na1185_6), .POUTY1(na1185_7), .POUTY2(na1185_8),
                      .IN1(na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1164_3), .CINY1(na1184_4), .CINY2(na1184_5), .PINX(na1164_6), .PINY1(na1184_7), .PINY2(na1184_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1186_1 ( .COUTX(na1186_3), .COUTY1(na1186_4), .COUTY2(na1186_5), .POUTX(na1186_6), .POUTY1(na1186_7), .POUTY2(na1186_8),
                      .IN1(~na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1165_3), .CINY1(na1185_4), .CINY2(na1185_5), .PINX(na1165_6), .PINY1(na1185_7), .PINY2(na1185_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1187_1 ( .COUTX(na1187_3), .COUTY1(na1187_4), .COUTY2(na1187_5), .POUTX(na1187_6), .POUTY1(na1187_7), .POUTY2(na1187_8),
                      .IN1(na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1166_3), .CINY1(na1186_4), .CINY2(na1186_5), .PINX(na1166_6), .PINY1(na1186_7), .PINY2(na1186_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1188_1 ( .COUTX(na1188_3), .COUTY1(na1188_4), .COUTY2(na1188_5), .POUTX(na1188_6), .POUTY1(na1188_7), .POUTY2(na1188_8),
                      .IN1(~na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1167_3), .CINY1(na1187_4), .CINY2(na1187_5), .PINX(na1167_6), .PINY1(na1187_7), .PINY2(na1187_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1189_1 ( .COUTX(na1189_3), .COUTY1(na1189_4), .COUTY2(na1189_5), .POUTX(na1189_6), .POUTY1(na1189_7), .POUTY2(na1189_8),
                      .IN1(na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1168_3), .CINY1(na1188_4), .CINY2(na1188_5), .PINX(na1168_6), .PINY1(na1188_7), .PINY2(na1188_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x28y58     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1190_1 ( .COUTX(na1190_3), .COUTY1(na1190_4), .COUTY2(na1190_5), .POUTX(na1190_6), .POUTY1(na1190_7), .POUTY2(na1190_8),
                      .IN1(~na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1169_3), .CINY1(na1189_4), .CINY2(na1189_5), .PINX(na1169_6), .PINY1(na1189_7), .PINY2(na1189_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x28y59     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1191_3 ( .COMP_OUT(na1191_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1191_4 ( .OUT(na1191_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1190_4), .PINX(1'b0), .PINY1(na1190_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1191_6 ( .COUTX(na1191_3), .POUTX(na1191_6), .CINX(1'b0), .CINY1(na1190_4), .CINY2(na1190_5), .PINX(1'b0), .PINY1(na1190_7),
                      .PINY2(na1190_8), .OUT1(1'b0), .OUT2(na1191_2), .COMP_OUT(na1191_3_i) );
// C_AND///AND/      x29y39     80'h00_0078_12_0000_0C88_FFF0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1192_1 ( .OUT(na1192_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1192_4 ( .OUT(na1192_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1192_6 ( .COUTY1(na1192_4), .POUTY1(na1192_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1192_1), .OUT2(na1192_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x29y40     80'h00_0018_04_2056_5888_0CCF
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1193_1 ( .OUT(na1193_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(na1172_3), .CINY1(na1192_4), .PINX(1'b0), .PINY1(na1192_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1193_3 ( .COMP_OUT(na1193_3_i), .COMB1(na1193_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1193_6 ( .COUTY1(na1193_4), .COUTY2(na1193_5), .POUTY1(na1193_7), .CINX(na1172_3), .CINY1(na1192_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1192_7), .PINY2(1'b0), .OUT1(na1193_1), .OUT2(1'b0), .COMP_OUT(na1193_3_i) );
// C_MULTFa//O_O2//      x29y41     80'h00_0018_13_A477_34A6_0CCC
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1194_1 ( .COUTX(na1194_3), .COUTY1(na1194_4), .COUTY2(na1194_5), .POUTY1(na1194_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1173_3), .CINY1(na1193_4),
                      .CINY2(na1193_5), .PINX(1'b0), .PINY1(na1193_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x29y42     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1195_1 ( .OUT(na1195_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1194_4), .PINX(1'b0), .PINY1(na1194_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1195_3 ( .COMP_OUT(na1195_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1195_4 ( .OUT(na1195_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1194_4), .PINX(1'b0), .PINY1(na1194_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1195_6 ( .COUTX(na1195_3), .COUTY1(na1195_4), .COUTY2(na1195_5), .POUTY1(na1195_7), .POUTY2(na1195_8), .CINX(1'b0), .CINY1(na1194_4),
                      .CINY2(na1194_5), .PINX(1'b0), .PINY1(na1194_7), .PINY2(1'b0), .OUT1(na1195_1), .OUT2(na1195_2), .COMP_OUT(na1195_3_i) );
// C_MULT///MULT/      x29y43     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1196_1 ( .COUTY1(na1196_4), .COUTY2(na1196_5), .POUTY1(na1196_7), .POUTY2(na1196_8), .IN1(na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1175_3),
                      .CINY1(na1195_4), .CINY2(na1195_5), .PINX(na1175_6), .PINY1(na1195_7), .PINY2(na1195_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y44     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1197_1 ( .COUTX(na1197_3), .COUTY1(na1197_4), .COUTY2(na1197_5), .POUTX(na1197_6), .POUTY1(na1197_7), .POUTY2(na1197_8),
                      .IN1(~na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1176_3), .CINY1(na1196_4), .CINY2(na1196_5), .PINX(na1176_6), .PINY1(na1196_7), .PINY2(na1196_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y45     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1198_1 ( .COUTX(na1198_3), .COUTY1(na1198_4), .COUTY2(na1198_5), .POUTX(na1198_6), .POUTY1(na1198_7), .POUTY2(na1198_8),
                      .IN1(na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1177_3), .CINY1(na1197_4), .CINY2(na1197_5), .PINX(na1177_6), .PINY1(na1197_7), .PINY2(na1197_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y46     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1199_1 ( .COUTX(na1199_3), .COUTY1(na1199_4), .COUTY2(na1199_5), .POUTX(na1199_6), .POUTY1(na1199_7), .POUTY2(na1199_8),
                      .IN1(~na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1178_3), .CINY1(na1198_4), .CINY2(na1198_5), .PINX(na1178_6), .PINY1(na1198_7), .PINY2(na1198_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y47     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1200_1 ( .COUTX(na1200_3), .COUTY1(na1200_4), .COUTY2(na1200_5), .POUTX(na1200_6), .POUTY1(na1200_7), .POUTY2(na1200_8),
                      .IN1(na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1179_3), .CINY1(na1199_4), .CINY2(na1199_5), .PINX(na1179_6), .PINY1(na1199_7), .PINY2(na1199_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y48     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1201_1 ( .COUTX(na1201_3), .COUTY1(na1201_4), .COUTY2(na1201_5), .POUTX(na1201_6), .POUTY1(na1201_7), .POUTY2(na1201_8),
                      .IN1(~na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1180_3), .CINY1(na1200_4), .CINY2(na1200_5), .PINX(na1180_6), .PINY1(na1200_7), .PINY2(na1200_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y49     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1202_1 ( .COUTX(na1202_3), .COUTY1(na1202_4), .COUTY2(na1202_5), .POUTX(na1202_6), .POUTY1(na1202_7), .POUTY2(na1202_8),
                      .IN1(na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1181_3), .CINY1(na1201_4), .CINY2(na1201_5), .PINX(na1181_6), .PINY1(na1201_7), .PINY2(na1201_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y50     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1203_1 ( .COUTX(na1203_3), .COUTY1(na1203_4), .COUTY2(na1203_5), .POUTX(na1203_6), .POUTY1(na1203_7), .POUTY2(na1203_8),
                      .IN1(~na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1182_3), .CINY1(na1202_4), .CINY2(na1202_5), .PINX(na1182_6), .PINY1(na1202_7), .PINY2(na1202_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y51     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1204_1 ( .COUTX(na1204_3), .COUTY1(na1204_4), .COUTY2(na1204_5), .POUTX(na1204_6), .POUTY1(na1204_7), .POUTY2(na1204_8),
                      .IN1(na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1183_3), .CINY1(na1203_4), .CINY2(na1203_5), .PINX(na1183_6), .PINY1(na1203_7), .PINY2(na1203_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y52     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1205_1 ( .COUTX(na1205_3), .COUTY1(na1205_4), .COUTY2(na1205_5), .POUTX(na1205_6), .POUTY1(na1205_7), .POUTY2(na1205_8),
                      .IN1(~na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1184_3), .CINY1(na1204_4), .CINY2(na1204_5), .PINX(na1184_6), .PINY1(na1204_7), .PINY2(na1204_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1206_1 ( .COUTX(na1206_3), .COUTY1(na1206_4), .COUTY2(na1206_5), .POUTX(na1206_6), .POUTY1(na1206_7), .POUTY2(na1206_8),
                      .IN1(na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1185_3), .CINY1(na1205_4), .CINY2(na1205_5), .PINX(na1185_6), .PINY1(na1205_7), .PINY2(na1205_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1207_1 ( .COUTX(na1207_3), .COUTY1(na1207_4), .COUTY2(na1207_5), .POUTX(na1207_6), .POUTY1(na1207_7), .POUTY2(na1207_8),
                      .IN1(~na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1186_3), .CINY1(na1206_4), .CINY2(na1206_5), .PINX(na1186_6), .PINY1(na1206_7), .PINY2(na1206_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1208_1 ( .COUTX(na1208_3), .COUTY1(na1208_4), .COUTY2(na1208_5), .POUTX(na1208_6), .POUTY1(na1208_7), .POUTY2(na1208_8),
                      .IN1(na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1187_3), .CINY1(na1207_4), .CINY2(na1207_5), .PINX(na1187_6), .PINY1(na1207_7), .PINY2(na1207_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1209_1 ( .COUTX(na1209_3), .COUTY1(na1209_4), .COUTY2(na1209_5), .POUTX(na1209_6), .POUTY1(na1209_7), .POUTY2(na1209_8),
                      .IN1(~na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1188_3), .CINY1(na1208_4), .CINY2(na1208_5), .PINX(na1188_6), .PINY1(na1208_7), .PINY2(na1208_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1210_1 ( .COUTX(na1210_3), .COUTY1(na1210_4), .COUTY2(na1210_5), .POUTX(na1210_6), .POUTY1(na1210_7), .POUTY2(na1210_8),
                      .IN1(na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1189_3), .CINY1(na1209_4), .CINY2(na1209_5), .PINX(na1189_6), .PINY1(na1209_7), .PINY2(na1209_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1211_1 ( .COUTX(na1211_3), .COUTY1(na1211_4), .COUTY2(na1211_5), .POUTX(na1211_6), .POUTY1(na1211_7), .POUTY2(na1211_8),
                      .IN1(~na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1190_3), .CINY1(na1210_4), .CINY2(na1210_5), .PINX(na1190_6), .PINY1(na1210_7), .PINY2(na1210_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x29y59     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1212_1 ( .COUTX(na1212_3), .COUTY1(na1212_4), .COUTY2(na1212_5), .POUTX(na1212_6), .POUTY1(na1212_7), .POUTY2(na1212_8),
                      .IN1(na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1191_3), .CINY1(na1211_4), .CINY2(na1211_5), .PINX(na1191_6), .PINY1(na1211_7), .PINY2(na1211_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x29y60     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1213_3 ( .COMP_OUT(na1213_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1213_4 ( .OUT(na1213_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1212_4), .PINX(1'b0), .PINY1(na1212_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1213_6 ( .COUTX(na1213_3), .POUTX(na1213_6), .CINX(1'b0), .CINY1(na1212_4), .CINY2(na1212_5), .PINX(1'b0), .PINY1(na1212_7),
                      .PINY2(na1212_8), .OUT1(1'b0), .OUT2(na1213_2), .COMP_OUT(na1213_3_i) );
// C_AND///AND/      x30y40     80'h00_0078_12_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1214_1 ( .OUT(na1214_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1214_4 ( .OUT(na1214_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1214_6 ( .COUTY1(na1214_4), .POUTY1(na1214_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1214_1), .OUT2(na1214_2), .COMP_OUT(1'b0) );
// C_OR//O_O1//      x30y41     80'h00_0018_04_2056_5EEE_0CC0
C_OR       #(.CPE_CFG (9'b0_0001_0110)) 
           _a1215_1 ( .OUT(na1215_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(na1194_3), .CINY1(na1214_4), .PINX(1'b0), .PINY1(na1214_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1215_3 ( .COMP_OUT(na1215_3_i), .COMB1(na1215_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1215_6 ( .COUTY1(na1215_4), .COUTY2(na1215_5), .POUTY1(na1215_7), .CINX(na1194_3), .CINY1(na1214_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1214_7), .PINY2(1'b0), .OUT1(na1215_1), .OUT2(1'b0), .COMP_OUT(na1215_3_i) );
// C_MULTFb//O_O2//      x30y42     80'h00_0018_13_A477_3EA6_0CCC
C_MULTFb   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1216_1 ( .COUTX(na1216_3), .COUTY1(na1216_4), .COUTY2(na1216_5), .POUTY1(na1216_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1195_3), .CINY1(na1215_4),
                      .CINY2(na1215_5), .PINX(1'b0), .PINY1(na1215_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_O2/AND/      x30y43     80'h00_0078_35_A471_3C88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1217_1 ( .OUT(na1217_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1216_4), .PINX(1'b0), .PINY1(na1216_7) );
C_O_O2     #(.CPE_CFG ()) 
           _a1217_3 ( .COMP_OUT(na1217_3_i), .COMB1(1'b0), .COMB2(na1217_2) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1217_4 ( .OUT(na1217_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1216_4), .PINX(1'b0), .PINY1(na1216_7) );
C_CPlines  #(.CPE_CFG (19'h3_5A47)) 
           _a1217_6 ( .COUTX(na1217_3), .COUTY1(na1217_4), .COUTY2(na1217_5), .POUTY1(na1217_7), .POUTY2(na1217_8), .CINX(1'b0), .CINY1(na1216_4),
                      .CINY2(na1216_5), .PINX(1'b0), .PINY1(na1216_7), .PINY2(1'b0), .OUT1(na1217_1), .OUT2(na1217_2), .COMP_OUT(na1217_3_i) );
// C_MULT///MULT/      x30y44     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1218_1 ( .COUTY1(na1218_4), .COUTY2(na1218_5), .POUTY1(na1218_7), .POUTY2(na1218_8), .IN1(~na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1197_3),
                      .CINY1(na1217_4), .CINY2(na1217_5), .PINX(na1197_6), .PINY1(na1217_7), .PINY2(na1217_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y45     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1219_1 ( .COUTX(na1219_3), .COUTY1(na1219_4), .COUTY2(na1219_5), .POUTX(na1219_6), .POUTY1(na1219_7), .POUTY2(na1219_8),
                      .IN1(na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1198_3), .CINY1(na1218_4), .CINY2(na1218_5), .PINX(na1198_6), .PINY1(na1218_7), .PINY2(na1218_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y46     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1220_1 ( .COUTX(na1220_3), .COUTY1(na1220_4), .COUTY2(na1220_5), .POUTX(na1220_6), .POUTY1(na1220_7), .POUTY2(na1220_8),
                      .IN1(~na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1199_3), .CINY1(na1219_4), .CINY2(na1219_5), .PINX(na1199_6), .PINY1(na1219_7), .PINY2(na1219_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y47     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1221_1 ( .COUTX(na1221_3), .COUTY1(na1221_4), .COUTY2(na1221_5), .POUTX(na1221_6), .POUTY1(na1221_7), .POUTY2(na1221_8),
                      .IN1(na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1200_3), .CINY1(na1220_4), .CINY2(na1220_5), .PINX(na1200_6), .PINY1(na1220_7), .PINY2(na1220_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y48     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1222_1 ( .COUTX(na1222_3), .COUTY1(na1222_4), .COUTY2(na1222_5), .POUTX(na1222_6), .POUTY1(na1222_7), .POUTY2(na1222_8),
                      .IN1(~na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1201_3), .CINY1(na1221_4), .CINY2(na1221_5), .PINX(na1201_6), .PINY1(na1221_7), .PINY2(na1221_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y49     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1223_1 ( .COUTX(na1223_3), .COUTY1(na1223_4), .COUTY2(na1223_5), .POUTX(na1223_6), .POUTY1(na1223_7), .POUTY2(na1223_8),
                      .IN1(na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1202_3), .CINY1(na1222_4), .CINY2(na1222_5), .PINX(na1202_6), .PINY1(na1222_7), .PINY2(na1222_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y50     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1224_1 ( .COUTX(na1224_3), .COUTY1(na1224_4), .COUTY2(na1224_5), .POUTX(na1224_6), .POUTY1(na1224_7), .POUTY2(na1224_8),
                      .IN1(~na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1203_3), .CINY1(na1223_4), .CINY2(na1223_5), .PINX(na1203_6), .PINY1(na1223_7), .PINY2(na1223_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y51     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1225_1 ( .COUTX(na1225_3), .COUTY1(na1225_4), .COUTY2(na1225_5), .POUTX(na1225_6), .POUTY1(na1225_7), .POUTY2(na1225_8),
                      .IN1(na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1204_3), .CINY1(na1224_4), .CINY2(na1224_5), .PINX(na1204_6), .PINY1(na1224_7), .PINY2(na1224_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y52     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1226_1 ( .COUTX(na1226_3), .COUTY1(na1226_4), .COUTY2(na1226_5), .POUTX(na1226_6), .POUTY1(na1226_7), .POUTY2(na1226_8),
                      .IN1(~na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1205_3), .CINY1(na1225_4), .CINY2(na1225_5), .PINX(na1205_6), .PINY1(na1225_7), .PINY2(na1225_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1227_1 ( .COUTX(na1227_3), .COUTY1(na1227_4), .COUTY2(na1227_5), .POUTX(na1227_6), .POUTY1(na1227_7), .POUTY2(na1227_8),
                      .IN1(na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1206_3), .CINY1(na1226_4), .CINY2(na1226_5), .PINX(na1206_6), .PINY1(na1226_7), .PINY2(na1226_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1228_1 ( .COUTX(na1228_3), .COUTY1(na1228_4), .COUTY2(na1228_5), .POUTX(na1228_6), .POUTY1(na1228_7), .POUTY2(na1228_8),
                      .IN1(~na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1207_3), .CINY1(na1227_4), .CINY2(na1227_5), .PINX(na1207_6), .PINY1(na1227_7), .PINY2(na1227_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1229_1 ( .COUTX(na1229_3), .COUTY1(na1229_4), .COUTY2(na1229_5), .POUTX(na1229_6), .POUTY1(na1229_7), .POUTY2(na1229_8),
                      .IN1(na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1208_3), .CINY1(na1228_4), .CINY2(na1228_5), .PINX(na1208_6), .PINY1(na1228_7), .PINY2(na1228_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1230_1 ( .COUTX(na1230_3), .COUTY1(na1230_4), .COUTY2(na1230_5), .POUTX(na1230_6), .POUTY1(na1230_7), .POUTY2(na1230_8),
                      .IN1(~na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1209_3), .CINY1(na1229_4), .CINY2(na1229_5), .PINX(na1209_6), .PINY1(na1229_7), .PINY2(na1229_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1231_1 ( .COUTX(na1231_3), .COUTY1(na1231_4), .COUTY2(na1231_5), .POUTX(na1231_6), .POUTY1(na1231_7), .POUTY2(na1231_8),
                      .IN1(na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1210_3), .CINY1(na1230_4), .CINY2(na1230_5), .PINX(na1210_6), .PINY1(na1230_7), .PINY2(na1230_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1232_1 ( .COUTX(na1232_3), .COUTY1(na1232_4), .COUTY2(na1232_5), .POUTX(na1232_6), .POUTY1(na1232_7), .POUTY2(na1232_8),
                      .IN1(~na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1211_3), .CINY1(na1231_4), .CINY2(na1231_5), .PINX(na1211_6), .PINY1(na1231_7), .PINY2(na1231_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1233_1 ( .COUTX(na1233_3), .COUTY1(na1233_4), .COUTY2(na1233_5), .POUTX(na1233_6), .POUTY1(na1233_7), .POUTY2(na1233_8),
                      .IN1(na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1212_3), .CINY1(na1232_4), .CINY2(na1232_5), .PINX(na1212_6), .PINY1(na1232_7), .PINY2(na1232_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x30y60     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1234_1 ( .COUTX(na1234_3), .COUTY1(na1234_4), .COUTY2(na1234_5), .POUTX(na1234_6), .POUTY1(na1234_7), .POUTY2(na1234_8),
                      .IN1(~na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1213_3), .CINY1(na1233_4), .CINY2(na1233_5), .PINX(na1213_6), .PINY1(na1233_7), .PINY2(na1233_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x30y61     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1235_3 ( .COMP_OUT(na1235_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1235_4 ( .OUT(na1235_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1234_4), .PINX(1'b0), .PINY1(na1234_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1235_6 ( .COUTX(na1235_3), .POUTX(na1235_6), .CINX(1'b0), .CINY1(na1234_4), .CINY2(na1234_5), .PINX(1'b0), .PINY1(na1234_7),
                      .PINY2(na1234_8), .OUT1(1'b0), .OUT2(na1235_2), .COMP_OUT(na1235_3_i) );
// C_AND///AND/      x31y41     80'h00_0078_12_0000_0C88_FFF0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1236_1 ( .OUT(na1236_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1236_4 ( .OUT(na1236_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1236_6 ( .COUTY1(na1236_4), .POUTY1(na1236_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1236_1), .OUT2(na1236_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x31y42     80'h00_0018_04_2056_5888_0CCF
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1237_1 ( .OUT(na1237_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(na1216_3), .CINY1(na1236_4), .PINX(1'b0), .PINY1(na1236_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1237_3 ( .COMP_OUT(na1237_3_i), .COMB1(na1237_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1237_6 ( .COUTY1(na1237_4), .COUTY2(na1237_5), .POUTY1(na1237_7), .CINX(na1216_3), .CINY1(na1236_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1236_7), .PINY2(1'b0), .OUT1(na1237_1), .OUT2(1'b0), .COMP_OUT(na1237_3_i) );
// C_MULTFa//O_O2//      x31y43     80'h00_0018_13_A477_34A6_0CCC
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1238_1 ( .COUTX(na1238_3), .COUTY1(na1238_4), .COUTY2(na1238_5), .POUTY1(na1238_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1217_3), .CINY1(na1237_4),
                      .CINY2(na1237_5), .PINX(1'b0), .PINY1(na1237_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x31y44     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1239_1 ( .OUT(na1239_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1238_4), .PINX(1'b0), .PINY1(na1238_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1239_3 ( .COMP_OUT(na1239_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1239_4 ( .OUT(na1239_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1238_4), .PINX(1'b0), .PINY1(na1238_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1239_6 ( .COUTX(na1239_3), .COUTY1(na1239_4), .COUTY2(na1239_5), .POUTY1(na1239_7), .POUTY2(na1239_8), .CINX(1'b0), .CINY1(na1238_4),
                      .CINY2(na1238_5), .PINX(1'b0), .PINY1(na1238_7), .PINY2(1'b0), .OUT1(na1239_1), .OUT2(na1239_2), .COMP_OUT(na1239_3_i) );
// C_MULT///MULT/      x31y45     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1240_1 ( .COUTY1(na1240_4), .COUTY2(na1240_5), .POUTY1(na1240_7), .POUTY2(na1240_8), .IN1(na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1219_3),
                      .CINY1(na1239_4), .CINY2(na1239_5), .PINX(na1219_6), .PINY1(na1239_7), .PINY2(na1239_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y46     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1241_1 ( .COUTX(na1241_3), .COUTY1(na1241_4), .COUTY2(na1241_5), .POUTX(na1241_6), .POUTY1(na1241_7), .POUTY2(na1241_8),
                      .IN1(~na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1220_3), .CINY1(na1240_4), .CINY2(na1240_5), .PINX(na1220_6), .PINY1(na1240_7), .PINY2(na1240_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y47     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1242_1 ( .COUTX(na1242_3), .COUTY1(na1242_4), .COUTY2(na1242_5), .POUTX(na1242_6), .POUTY1(na1242_7), .POUTY2(na1242_8),
                      .IN1(na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1221_3), .CINY1(na1241_4), .CINY2(na1241_5), .PINX(na1221_6), .PINY1(na1241_7), .PINY2(na1241_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y48     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1243_1 ( .COUTX(na1243_3), .COUTY1(na1243_4), .COUTY2(na1243_5), .POUTX(na1243_6), .POUTY1(na1243_7), .POUTY2(na1243_8),
                      .IN1(~na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1222_3), .CINY1(na1242_4), .CINY2(na1242_5), .PINX(na1222_6), .PINY1(na1242_7), .PINY2(na1242_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y49     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1244_1 ( .COUTX(na1244_3), .COUTY1(na1244_4), .COUTY2(na1244_5), .POUTX(na1244_6), .POUTY1(na1244_7), .POUTY2(na1244_8),
                      .IN1(na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1223_3), .CINY1(na1243_4), .CINY2(na1243_5), .PINX(na1223_6), .PINY1(na1243_7), .PINY2(na1243_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y50     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1245_1 ( .COUTX(na1245_3), .COUTY1(na1245_4), .COUTY2(na1245_5), .POUTX(na1245_6), .POUTY1(na1245_7), .POUTY2(na1245_8),
                      .IN1(~na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1224_3), .CINY1(na1244_4), .CINY2(na1244_5), .PINX(na1224_6), .PINY1(na1244_7), .PINY2(na1244_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y51     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1246_1 ( .COUTX(na1246_3), .COUTY1(na1246_4), .COUTY2(na1246_5), .POUTX(na1246_6), .POUTY1(na1246_7), .POUTY2(na1246_8),
                      .IN1(na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1225_3), .CINY1(na1245_4), .CINY2(na1245_5), .PINX(na1225_6), .PINY1(na1245_7), .PINY2(na1245_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y52     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1247_1 ( .COUTX(na1247_3), .COUTY1(na1247_4), .COUTY2(na1247_5), .POUTX(na1247_6), .POUTY1(na1247_7), .POUTY2(na1247_8),
                      .IN1(~na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1226_3), .CINY1(na1246_4), .CINY2(na1246_5), .PINX(na1226_6), .PINY1(na1246_7), .PINY2(na1246_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1248_1 ( .COUTX(na1248_3), .COUTY1(na1248_4), .COUTY2(na1248_5), .POUTX(na1248_6), .POUTY1(na1248_7), .POUTY2(na1248_8),
                      .IN1(na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1227_3), .CINY1(na1247_4), .CINY2(na1247_5), .PINX(na1227_6), .PINY1(na1247_7), .PINY2(na1247_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1249_1 ( .COUTX(na1249_3), .COUTY1(na1249_4), .COUTY2(na1249_5), .POUTX(na1249_6), .POUTY1(na1249_7), .POUTY2(na1249_8),
                      .IN1(~na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1228_3), .CINY1(na1248_4), .CINY2(na1248_5), .PINX(na1228_6), .PINY1(na1248_7), .PINY2(na1248_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1250_1 ( .COUTX(na1250_3), .COUTY1(na1250_4), .COUTY2(na1250_5), .POUTX(na1250_6), .POUTY1(na1250_7), .POUTY2(na1250_8),
                      .IN1(na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1229_3), .CINY1(na1249_4), .CINY2(na1249_5), .PINX(na1229_6), .PINY1(na1249_7), .PINY2(na1249_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1251_1 ( .COUTX(na1251_3), .COUTY1(na1251_4), .COUTY2(na1251_5), .POUTX(na1251_6), .POUTY1(na1251_7), .POUTY2(na1251_8),
                      .IN1(~na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1230_3), .CINY1(na1250_4), .CINY2(na1250_5), .PINX(na1230_6), .PINY1(na1250_7), .PINY2(na1250_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1252_1 ( .COUTX(na1252_3), .COUTY1(na1252_4), .COUTY2(na1252_5), .POUTX(na1252_6), .POUTY1(na1252_7), .POUTY2(na1252_8),
                      .IN1(na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1231_3), .CINY1(na1251_4), .CINY2(na1251_5), .PINX(na1231_6), .PINY1(na1251_7), .PINY2(na1251_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1253_1 ( .COUTX(na1253_3), .COUTY1(na1253_4), .COUTY2(na1253_5), .POUTX(na1253_6), .POUTY1(na1253_7), .POUTY2(na1253_8),
                      .IN1(~na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1232_3), .CINY1(na1252_4), .CINY2(na1252_5), .PINX(na1232_6), .PINY1(na1252_7), .PINY2(na1252_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1254_1 ( .COUTX(na1254_3), .COUTY1(na1254_4), .COUTY2(na1254_5), .POUTX(na1254_6), .POUTY1(na1254_7), .POUTY2(na1254_8),
                      .IN1(na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1233_3), .CINY1(na1253_4), .CINY2(na1253_5), .PINX(na1233_6), .PINY1(na1253_7), .PINY2(na1253_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1255_1 ( .COUTX(na1255_3), .COUTY1(na1255_4), .COUTY2(na1255_5), .POUTX(na1255_6), .POUTY1(na1255_7), .POUTY2(na1255_8),
                      .IN1(~na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1234_3), .CINY1(na1254_4), .CINY2(na1254_5), .PINX(na1234_6), .PINY1(na1254_7), .PINY2(na1254_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x31y61     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1256_1 ( .COUTX(na1256_3), .COUTY1(na1256_4), .COUTY2(na1256_5), .POUTX(na1256_6), .POUTY1(na1256_7), .POUTY2(na1256_8),
                      .IN1(na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1235_3), .CINY1(na1255_4), .CINY2(na1255_5), .PINX(na1235_6), .PINY1(na1255_7), .PINY2(na1255_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x31y62     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1257_3 ( .COMP_OUT(na1257_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1257_4 ( .OUT(na1257_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1256_4), .PINX(1'b0), .PINY1(na1256_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1257_6 ( .COUTX(na1257_3), .POUTX(na1257_6), .CINX(1'b0), .CINY1(na1256_4), .CINY2(na1256_5), .PINX(1'b0), .PINY1(na1256_7),
                      .PINY2(na1256_8), .OUT1(1'b0), .OUT2(na1257_2), .COMP_OUT(na1257_3_i) );
// C_AND///AND/      x32y42     80'h00_0078_12_0000_0C88_F0F0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1258_1 ( .OUT(na1258_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1258_4 ( .OUT(na1258_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1258_6 ( .COUTY1(na1258_4), .POUTY1(na1258_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1258_1), .OUT2(na1258_2), .COMP_OUT(1'b0) );
// C_OR//O_O1//      x32y43     80'h00_0018_04_2056_5EEE_0CC0
C_OR       #(.CPE_CFG (9'b0_0001_0110)) 
           _a1259_1 ( .OUT(na1259_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(na1238_3), .CINY1(na1258_4), .PINX(1'b0), .PINY1(na1258_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1259_3 ( .COMP_OUT(na1259_3_i), .COMB1(na1259_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1259_6 ( .COUTY1(na1259_4), .COUTY2(na1259_5), .POUTY1(na1259_7), .CINX(na1238_3), .CINY1(na1258_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1258_7), .PINY2(1'b0), .OUT1(na1259_1), .OUT2(1'b0), .COMP_OUT(na1259_3_i) );
// C_MULTFb//O_O2//      x32y44     80'h00_0018_13_A477_3EA6_0CCC
C_MULTFb   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1260_1 ( .COUTX(na1260_3), .COUTY1(na1260_4), .COUTY2(na1260_5), .POUTY1(na1260_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1239_3), .CINY1(na1259_4),
                      .CINY2(na1259_5), .PINX(1'b0), .PINY1(na1259_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_O2/AND/      x32y45     80'h00_0078_35_A471_3C88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1261_1 ( .OUT(na1261_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1260_4), .PINX(1'b0), .PINY1(na1260_7) );
C_O_O2     #(.CPE_CFG ()) 
           _a1261_3 ( .COMP_OUT(na1261_3_i), .COMB1(1'b0), .COMB2(na1261_2) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1261_4 ( .OUT(na1261_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1260_4), .PINX(1'b0), .PINY1(na1260_7) );
C_CPlines  #(.CPE_CFG (19'h3_5A47)) 
           _a1261_6 ( .COUTX(na1261_3), .COUTY1(na1261_4), .COUTY2(na1261_5), .POUTY1(na1261_7), .POUTY2(na1261_8), .CINX(1'b0), .CINY1(na1260_4),
                      .CINY2(na1260_5), .PINX(1'b0), .PINY1(na1260_7), .PINY2(1'b0), .OUT1(na1261_1), .OUT2(na1261_2), .COMP_OUT(na1261_3_i) );
// C_MULT///MULT/      x32y46     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1262_1 ( .COUTY1(na1262_4), .COUTY2(na1262_5), .POUTY1(na1262_7), .POUTY2(na1262_8), .IN1(~na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1241_3),
                      .CINY1(na1261_4), .CINY2(na1261_5), .PINX(na1241_6), .PINY1(na1261_7), .PINY2(na1261_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y47     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1263_1 ( .COUTX(na1263_3), .COUTY1(na1263_4), .COUTY2(na1263_5), .POUTX(na1263_6), .POUTY1(na1263_7), .POUTY2(na1263_8),
                      .IN1(na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1242_3), .CINY1(na1262_4), .CINY2(na1262_5), .PINX(na1242_6), .PINY1(na1262_7), .PINY2(na1262_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y48     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1264_1 ( .COUTX(na1264_3), .COUTY1(na1264_4), .COUTY2(na1264_5), .POUTX(na1264_6), .POUTY1(na1264_7), .POUTY2(na1264_8),
                      .IN1(~na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1243_3), .CINY1(na1263_4), .CINY2(na1263_5), .PINX(na1243_6), .PINY1(na1263_7), .PINY2(na1263_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y49     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1265_1 ( .COUTX(na1265_3), .COUTY1(na1265_4), .COUTY2(na1265_5), .POUTX(na1265_6), .POUTY1(na1265_7), .POUTY2(na1265_8),
                      .IN1(na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1244_3), .CINY1(na1264_4), .CINY2(na1264_5), .PINX(na1244_6), .PINY1(na1264_7), .PINY2(na1264_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y50     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1266_1 ( .COUTX(na1266_3), .COUTY1(na1266_4), .COUTY2(na1266_5), .POUTX(na1266_6), .POUTY1(na1266_7), .POUTY2(na1266_8),
                      .IN1(~na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1245_3), .CINY1(na1265_4), .CINY2(na1265_5), .PINX(na1245_6), .PINY1(na1265_7), .PINY2(na1265_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y51     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1267_1 ( .COUTX(na1267_3), .COUTY1(na1267_4), .COUTY2(na1267_5), .POUTX(na1267_6), .POUTY1(na1267_7), .POUTY2(na1267_8),
                      .IN1(na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1246_3), .CINY1(na1266_4), .CINY2(na1266_5), .PINX(na1246_6), .PINY1(na1266_7), .PINY2(na1266_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y52     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1268_1 ( .COUTX(na1268_3), .COUTY1(na1268_4), .COUTY2(na1268_5), .POUTX(na1268_6), .POUTY1(na1268_7), .POUTY2(na1268_8),
                      .IN1(~na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1247_3), .CINY1(na1267_4), .CINY2(na1267_5), .PINX(na1247_6), .PINY1(na1267_7), .PINY2(na1267_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1269_1 ( .COUTX(na1269_3), .COUTY1(na1269_4), .COUTY2(na1269_5), .POUTX(na1269_6), .POUTY1(na1269_7), .POUTY2(na1269_8),
                      .IN1(na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1248_3), .CINY1(na1268_4), .CINY2(na1268_5), .PINX(na1248_6), .PINY1(na1268_7), .PINY2(na1268_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1270_1 ( .COUTX(na1270_3), .COUTY1(na1270_4), .COUTY2(na1270_5), .POUTX(na1270_6), .POUTY1(na1270_7), .POUTY2(na1270_8),
                      .IN1(~na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1249_3), .CINY1(na1269_4), .CINY2(na1269_5), .PINX(na1249_6), .PINY1(na1269_7), .PINY2(na1269_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1271_1 ( .COUTX(na1271_3), .COUTY1(na1271_4), .COUTY2(na1271_5), .POUTX(na1271_6), .POUTY1(na1271_7), .POUTY2(na1271_8),
                      .IN1(na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1250_3), .CINY1(na1270_4), .CINY2(na1270_5), .PINX(na1250_6), .PINY1(na1270_7), .PINY2(na1270_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1272_1 ( .COUTX(na1272_3), .COUTY1(na1272_4), .COUTY2(na1272_5), .POUTX(na1272_6), .POUTY1(na1272_7), .POUTY2(na1272_8),
                      .IN1(~na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1251_3), .CINY1(na1271_4), .CINY2(na1271_5), .PINX(na1251_6), .PINY1(na1271_7), .PINY2(na1271_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1273_1 ( .COUTX(na1273_3), .COUTY1(na1273_4), .COUTY2(na1273_5), .POUTX(na1273_6), .POUTY1(na1273_7), .POUTY2(na1273_8),
                      .IN1(na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1252_3), .CINY1(na1272_4), .CINY2(na1272_5), .PINX(na1252_6), .PINY1(na1272_7), .PINY2(na1272_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1274_1 ( .COUTX(na1274_3), .COUTY1(na1274_4), .COUTY2(na1274_5), .POUTX(na1274_6), .POUTY1(na1274_7), .POUTY2(na1274_8),
                      .IN1(~na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1253_3), .CINY1(na1273_4), .CINY2(na1273_5), .PINX(na1253_6), .PINY1(na1273_7), .PINY2(na1273_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1275_1 ( .COUTX(na1275_3), .COUTY1(na1275_4), .COUTY2(na1275_5), .POUTX(na1275_6), .POUTY1(na1275_7), .POUTY2(na1275_8),
                      .IN1(na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1254_3), .CINY1(na1274_4), .CINY2(na1274_5), .PINX(na1254_6), .PINY1(na1274_7), .PINY2(na1274_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1276_1 ( .COUTX(na1276_3), .COUTY1(na1276_4), .COUTY2(na1276_5), .POUTX(na1276_6), .POUTY1(na1276_7), .POUTY2(na1276_8),
                      .IN1(~na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1255_3), .CINY1(na1275_4), .CINY2(na1275_5), .PINX(na1255_6), .PINY1(na1275_7), .PINY2(na1275_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y61     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1277_1 ( .COUTX(na1277_3), .COUTY1(na1277_4), .COUTY2(na1277_5), .POUTX(na1277_6), .POUTY1(na1277_7), .POUTY2(na1277_8),
                      .IN1(na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1256_3), .CINY1(na1276_4), .CINY2(na1276_5), .PINX(na1256_6), .PINY1(na1276_7), .PINY2(na1276_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x32y62     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1278_1 ( .COUTX(na1278_3), .COUTY1(na1278_4), .COUTY2(na1278_5), .POUTX(na1278_6), .POUTY1(na1278_7), .POUTY2(na1278_8),
                      .IN1(~na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1257_3), .CINY1(na1277_4), .CINY2(na1277_5), .PINX(na1257_6), .PINY1(na1277_7), .PINY2(na1277_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x32y63     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1279_3 ( .COMP_OUT(na1279_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1279_4 ( .OUT(na1279_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1278_4), .PINX(1'b0), .PINY1(na1278_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1279_6 ( .COUTX(na1279_3), .POUTX(na1279_6), .CINX(1'b0), .CINY1(na1278_4), .CINY2(na1278_5), .PINX(1'b0), .PINY1(na1278_7),
                      .PINY2(na1278_8), .OUT1(1'b0), .OUT2(na1279_2), .COMP_OUT(na1279_3_i) );
// C_AND///AND/      x33y43     80'h00_0078_12_0000_0C88_FFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1280_1 ( .OUT(na1280_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1280_4 ( .OUT(na1280_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1280_6 ( .COUTY1(na1280_4), .POUTY1(na1280_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1280_1), .OUT2(na1280_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x33y44     80'h00_0018_04_2056_5888_0CCF
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1281_1 ( .OUT(na1281_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(na1260_3), .CINY1(na1280_4), .PINX(1'b0), .PINY1(na1280_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1281_3 ( .COMP_OUT(na1281_3_i), .COMB1(na1281_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1281_6 ( .COUTY1(na1281_4), .COUTY2(na1281_5), .POUTY1(na1281_7), .CINX(na1260_3), .CINY1(na1280_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1280_7), .PINY2(1'b0), .OUT1(na1281_1), .OUT2(1'b0), .COMP_OUT(na1281_3_i) );
// C_MULTFa//O_O2//      x33y45     80'h00_0018_13_A477_34A6_0CCC
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1282_1 ( .COUTX(na1282_3), .COUTY1(na1282_4), .COUTY2(na1282_5), .POUTY1(na1282_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1261_3), .CINY1(na1281_4),
                      .CINY2(na1281_5), .PINX(1'b0), .PINY1(na1281_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x33y46     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1283_1 ( .OUT(na1283_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1282_4), .PINX(1'b0), .PINY1(na1282_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1283_3 ( .COMP_OUT(na1283_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1283_4 ( .OUT(na1283_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1282_4), .PINX(1'b0), .PINY1(na1282_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1283_6 ( .COUTX(na1283_3), .COUTY1(na1283_4), .COUTY2(na1283_5), .POUTY1(na1283_7), .POUTY2(na1283_8), .CINX(1'b0), .CINY1(na1282_4),
                      .CINY2(na1282_5), .PINX(1'b0), .PINY1(na1282_7), .PINY2(1'b0), .OUT1(na1283_1), .OUT2(na1283_2), .COMP_OUT(na1283_3_i) );
// C_MULT///MULT/      x33y47     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1284_1 ( .COUTY1(na1284_4), .COUTY2(na1284_5), .POUTY1(na1284_7), .POUTY2(na1284_8), .IN1(na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1263_3),
                      .CINY1(na1283_4), .CINY2(na1283_5), .PINX(na1263_6), .PINY1(na1283_7), .PINY2(na1283_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y48     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1285_1 ( .COUTX(na1285_3), .COUTY1(na1285_4), .COUTY2(na1285_5), .POUTX(na1285_6), .POUTY1(na1285_7), .POUTY2(na1285_8),
                      .IN1(~na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1264_3), .CINY1(na1284_4), .CINY2(na1284_5), .PINX(na1264_6), .PINY1(na1284_7), .PINY2(na1284_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y49     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1286_1 ( .COUTX(na1286_3), .COUTY1(na1286_4), .COUTY2(na1286_5), .POUTX(na1286_6), .POUTY1(na1286_7), .POUTY2(na1286_8),
                      .IN1(na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1265_3), .CINY1(na1285_4), .CINY2(na1285_5), .PINX(na1265_6), .PINY1(na1285_7), .PINY2(na1285_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y50     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1287_1 ( .COUTX(na1287_3), .COUTY1(na1287_4), .COUTY2(na1287_5), .POUTX(na1287_6), .POUTY1(na1287_7), .POUTY2(na1287_8),
                      .IN1(~na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1266_3), .CINY1(na1286_4), .CINY2(na1286_5), .PINX(na1266_6), .PINY1(na1286_7), .PINY2(na1286_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y51     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1288_1 ( .COUTX(na1288_3), .COUTY1(na1288_4), .COUTY2(na1288_5), .POUTX(na1288_6), .POUTY1(na1288_7), .POUTY2(na1288_8),
                      .IN1(na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1267_3), .CINY1(na1287_4), .CINY2(na1287_5), .PINX(na1267_6), .PINY1(na1287_7), .PINY2(na1287_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y52     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1289_1 ( .COUTX(na1289_3), .COUTY1(na1289_4), .COUTY2(na1289_5), .POUTX(na1289_6), .POUTY1(na1289_7), .POUTY2(na1289_8),
                      .IN1(~na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1268_3), .CINY1(na1288_4), .CINY2(na1288_5), .PINX(na1268_6), .PINY1(na1288_7), .PINY2(na1288_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1290_1 ( .COUTX(na1290_3), .COUTY1(na1290_4), .COUTY2(na1290_5), .POUTX(na1290_6), .POUTY1(na1290_7), .POUTY2(na1290_8),
                      .IN1(na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1269_3), .CINY1(na1289_4), .CINY2(na1289_5), .PINX(na1269_6), .PINY1(na1289_7), .PINY2(na1289_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1291_1 ( .COUTX(na1291_3), .COUTY1(na1291_4), .COUTY2(na1291_5), .POUTX(na1291_6), .POUTY1(na1291_7), .POUTY2(na1291_8),
                      .IN1(~na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1270_3), .CINY1(na1290_4), .CINY2(na1290_5), .PINX(na1270_6), .PINY1(na1290_7), .PINY2(na1290_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1292_1 ( .COUTX(na1292_3), .COUTY1(na1292_4), .COUTY2(na1292_5), .POUTX(na1292_6), .POUTY1(na1292_7), .POUTY2(na1292_8),
                      .IN1(na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1271_3), .CINY1(na1291_4), .CINY2(na1291_5), .PINX(na1271_6), .PINY1(na1291_7), .PINY2(na1291_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1293_1 ( .COUTX(na1293_3), .COUTY1(na1293_4), .COUTY2(na1293_5), .POUTX(na1293_6), .POUTY1(na1293_7), .POUTY2(na1293_8),
                      .IN1(~na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1272_3), .CINY1(na1292_4), .CINY2(na1292_5), .PINX(na1272_6), .PINY1(na1292_7), .PINY2(na1292_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1294_1 ( .COUTX(na1294_3), .COUTY1(na1294_4), .COUTY2(na1294_5), .POUTX(na1294_6), .POUTY1(na1294_7), .POUTY2(na1294_8),
                      .IN1(na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1273_3), .CINY1(na1293_4), .CINY2(na1293_5), .PINX(na1273_6), .PINY1(na1293_7), .PINY2(na1293_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1295_1 ( .COUTX(na1295_3), .COUTY1(na1295_4), .COUTY2(na1295_5), .POUTX(na1295_6), .POUTY1(na1295_7), .POUTY2(na1295_8),
                      .IN1(~na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1274_3), .CINY1(na1294_4), .CINY2(na1294_5), .PINX(na1274_6), .PINY1(na1294_7), .PINY2(na1294_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1296_1 ( .COUTX(na1296_3), .COUTY1(na1296_4), .COUTY2(na1296_5), .POUTX(na1296_6), .POUTY1(na1296_7), .POUTY2(na1296_8),
                      .IN1(na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1275_3), .CINY1(na1295_4), .CINY2(na1295_5), .PINX(na1275_6), .PINY1(na1295_7), .PINY2(na1295_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1297_1 ( .COUTX(na1297_3), .COUTY1(na1297_4), .COUTY2(na1297_5), .POUTX(na1297_6), .POUTY1(na1297_7), .POUTY2(na1297_8),
                      .IN1(~na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1276_3), .CINY1(na1296_4), .CINY2(na1296_5), .PINX(na1276_6), .PINY1(na1296_7), .PINY2(na1296_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y61     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1298_1 ( .COUTX(na1298_3), .COUTY1(na1298_4), .COUTY2(na1298_5), .POUTX(na1298_6), .POUTY1(na1298_7), .POUTY2(na1298_8),
                      .IN1(na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1277_3), .CINY1(na1297_4), .CINY2(na1297_5), .PINX(na1277_6), .PINY1(na1297_7), .PINY2(na1297_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y62     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1299_1 ( .COUTX(na1299_3), .COUTY1(na1299_4), .COUTY2(na1299_5), .POUTX(na1299_6), .POUTY1(na1299_7), .POUTY2(na1299_8),
                      .IN1(~na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1278_3), .CINY1(na1298_4), .CINY2(na1298_5), .PINX(na1278_6), .PINY1(na1298_7), .PINY2(na1298_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x33y63     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1300_1 ( .COUTX(na1300_3), .COUTY1(na1300_4), .COUTY2(na1300_5), .POUTX(na1300_6), .POUTY1(na1300_7), .POUTY2(na1300_8),
                      .IN1(na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1279_3), .CINY1(na1299_4), .CINY2(na1299_5), .PINX(na1279_6), .PINY1(na1299_7), .PINY2(na1299_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x33y64     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1301_3 ( .COMP_OUT(na1301_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1301_4 ( .OUT(na1301_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1300_4), .PINX(1'b0), .PINY1(na1300_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1301_6 ( .COUTX(na1301_3), .POUTX(na1301_6), .CINX(1'b0), .CINY1(na1300_4), .CINY2(na1300_5), .PINX(1'b0), .PINY1(na1300_7),
                      .PINY2(na1300_8), .OUT1(1'b0), .OUT2(na1301_2), .COMP_OUT(na1301_3_i) );
// C_AND///AND/      x34y44     80'h00_0078_12_0000_0C88_F0F0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1302_1 ( .OUT(na1302_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1302_4 ( .OUT(na1302_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1302_6 ( .COUTY1(na1302_4), .POUTY1(na1302_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1302_1), .OUT2(na1302_2), .COMP_OUT(1'b0) );
// C_OR//O_O1//      x34y45     80'h00_0018_04_2056_5EEE_0CC0
C_OR       #(.CPE_CFG (9'b0_0001_0110)) 
           _a1303_1 ( .OUT(na1303_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(na1282_3), .CINY1(na1302_4), .PINX(1'b0), .PINY1(na1302_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1303_3 ( .COMP_OUT(na1303_3_i), .COMB1(na1303_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1303_6 ( .COUTY1(na1303_4), .COUTY2(na1303_5), .POUTY1(na1303_7), .CINX(na1282_3), .CINY1(na1302_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1302_7), .PINY2(1'b0), .OUT1(na1303_1), .OUT2(1'b0), .COMP_OUT(na1303_3_i) );
// C_MULTFb//O_O2//      x34y46     80'h00_0018_13_A477_3EA6_0CCC
C_MULTFb   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1304_1 ( .COUTX(na1304_3), .COUTY1(na1304_4), .COUTY2(na1304_5), .POUTY1(na1304_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1283_3), .CINY1(na1303_4),
                      .CINY2(na1303_5), .PINX(1'b0), .PINY1(na1303_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_O2/AND/      x34y47     80'h00_0078_35_A471_3C88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1305_1 ( .OUT(na1305_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1304_4), .PINX(1'b0), .PINY1(na1304_7) );
C_O_O2     #(.CPE_CFG ()) 
           _a1305_3 ( .COMP_OUT(na1305_3_i), .COMB1(1'b0), .COMB2(na1305_2) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1305_4 ( .OUT(na1305_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1304_4), .PINX(1'b0), .PINY1(na1304_7) );
C_CPlines  #(.CPE_CFG (19'h3_5A47)) 
           _a1305_6 ( .COUTX(na1305_3), .COUTY1(na1305_4), .COUTY2(na1305_5), .POUTY1(na1305_7), .POUTY2(na1305_8), .CINX(1'b0), .CINY1(na1304_4),
                      .CINY2(na1304_5), .PINX(1'b0), .PINY1(na1304_7), .PINY2(1'b0), .OUT1(na1305_1), .OUT2(na1305_2), .COMP_OUT(na1305_3_i) );
// C_MULT///MULT/      x34y48     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1306_1 ( .COUTY1(na1306_4), .COUTY2(na1306_5), .POUTY1(na1306_7), .POUTY2(na1306_8), .IN1(~na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1285_3),
                      .CINY1(na1305_4), .CINY2(na1305_5), .PINX(na1285_6), .PINY1(na1305_7), .PINY2(na1305_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y49     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1307_1 ( .COUTX(na1307_3), .COUTY1(na1307_4), .COUTY2(na1307_5), .POUTX(na1307_6), .POUTY1(na1307_7), .POUTY2(na1307_8),
                      .IN1(na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1286_3), .CINY1(na1306_4), .CINY2(na1306_5), .PINX(na1286_6), .PINY1(na1306_7), .PINY2(na1306_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y50     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1308_1 ( .COUTX(na1308_3), .COUTY1(na1308_4), .COUTY2(na1308_5), .POUTX(na1308_6), .POUTY1(na1308_7), .POUTY2(na1308_8),
                      .IN1(~na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1287_3), .CINY1(na1307_4), .CINY2(na1307_5), .PINX(na1287_6), .PINY1(na1307_7), .PINY2(na1307_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y51     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1309_1 ( .COUTX(na1309_3), .COUTY1(na1309_4), .COUTY2(na1309_5), .POUTX(na1309_6), .POUTY1(na1309_7), .POUTY2(na1309_8),
                      .IN1(na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1288_3), .CINY1(na1308_4), .CINY2(na1308_5), .PINX(na1288_6), .PINY1(na1308_7), .PINY2(na1308_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y52     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1310_1 ( .COUTX(na1310_3), .COUTY1(na1310_4), .COUTY2(na1310_5), .POUTX(na1310_6), .POUTY1(na1310_7), .POUTY2(na1310_8),
                      .IN1(~na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1289_3), .CINY1(na1309_4), .CINY2(na1309_5), .PINX(na1289_6), .PINY1(na1309_7), .PINY2(na1309_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1311_1 ( .COUTX(na1311_3), .COUTY1(na1311_4), .COUTY2(na1311_5), .POUTX(na1311_6), .POUTY1(na1311_7), .POUTY2(na1311_8),
                      .IN1(na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1290_3), .CINY1(na1310_4), .CINY2(na1310_5), .PINX(na1290_6), .PINY1(na1310_7), .PINY2(na1310_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1312_1 ( .COUTX(na1312_3), .COUTY1(na1312_4), .COUTY2(na1312_5), .POUTX(na1312_6), .POUTY1(na1312_7), .POUTY2(na1312_8),
                      .IN1(~na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1291_3), .CINY1(na1311_4), .CINY2(na1311_5), .PINX(na1291_6), .PINY1(na1311_7), .PINY2(na1311_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1313_1 ( .COUTX(na1313_3), .COUTY1(na1313_4), .COUTY2(na1313_5), .POUTX(na1313_6), .POUTY1(na1313_7), .POUTY2(na1313_8),
                      .IN1(na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1292_3), .CINY1(na1312_4), .CINY2(na1312_5), .PINX(na1292_6), .PINY1(na1312_7), .PINY2(na1312_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1314_1 ( .COUTX(na1314_3), .COUTY1(na1314_4), .COUTY2(na1314_5), .POUTX(na1314_6), .POUTY1(na1314_7), .POUTY2(na1314_8),
                      .IN1(~na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1293_3), .CINY1(na1313_4), .CINY2(na1313_5), .PINX(na1293_6), .PINY1(na1313_7), .PINY2(na1313_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1315_1 ( .COUTX(na1315_3), .COUTY1(na1315_4), .COUTY2(na1315_5), .POUTX(na1315_6), .POUTY1(na1315_7), .POUTY2(na1315_8),
                      .IN1(na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1294_3), .CINY1(na1314_4), .CINY2(na1314_5), .PINX(na1294_6), .PINY1(na1314_7), .PINY2(na1314_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1316_1 ( .COUTX(na1316_3), .COUTY1(na1316_4), .COUTY2(na1316_5), .POUTX(na1316_6), .POUTY1(na1316_7), .POUTY2(na1316_8),
                      .IN1(~na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1295_3), .CINY1(na1315_4), .CINY2(na1315_5), .PINX(na1295_6), .PINY1(na1315_7), .PINY2(na1315_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1317_1 ( .COUTX(na1317_3), .COUTY1(na1317_4), .COUTY2(na1317_5), .POUTX(na1317_6), .POUTY1(na1317_7), .POUTY2(na1317_8),
                      .IN1(na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1296_3), .CINY1(na1316_4), .CINY2(na1316_5), .PINX(na1296_6), .PINY1(na1316_7), .PINY2(na1316_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1318_1 ( .COUTX(na1318_3), .COUTY1(na1318_4), .COUTY2(na1318_5), .POUTX(na1318_6), .POUTY1(na1318_7), .POUTY2(na1318_8),
                      .IN1(~na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1297_3), .CINY1(na1317_4), .CINY2(na1317_5), .PINX(na1297_6), .PINY1(na1317_7), .PINY2(na1317_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y61     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1319_1 ( .COUTX(na1319_3), .COUTY1(na1319_4), .COUTY2(na1319_5), .POUTX(na1319_6), .POUTY1(na1319_7), .POUTY2(na1319_8),
                      .IN1(na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1298_3), .CINY1(na1318_4), .CINY2(na1318_5), .PINX(na1298_6), .PINY1(na1318_7), .PINY2(na1318_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y62     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1320_1 ( .COUTX(na1320_3), .COUTY1(na1320_4), .COUTY2(na1320_5), .POUTX(na1320_6), .POUTY1(na1320_7), .POUTY2(na1320_8),
                      .IN1(~na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1299_3), .CINY1(na1319_4), .CINY2(na1319_5), .PINX(na1299_6), .PINY1(na1319_7), .PINY2(na1319_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y63     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1321_1 ( .COUTX(na1321_3), .COUTY1(na1321_4), .COUTY2(na1321_5), .POUTX(na1321_6), .POUTY1(na1321_7), .POUTY2(na1321_8),
                      .IN1(na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1300_3), .CINY1(na1320_4), .CINY2(na1320_5), .PINX(na1300_6), .PINY1(na1320_7), .PINY2(na1320_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x34y64     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1322_1 ( .COUTX(na1322_3), .COUTY1(na1322_4), .COUTY2(na1322_5), .POUTX(na1322_6), .POUTY1(na1322_7), .POUTY2(na1322_8),
                      .IN1(~na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1301_3), .CINY1(na1321_4), .CINY2(na1321_5), .PINX(na1301_6), .PINY1(na1321_7), .PINY2(na1321_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x34y65     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1323_3 ( .COMP_OUT(na1323_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1323_4 ( .OUT(na1323_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1322_4), .PINX(1'b0), .PINY1(na1322_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1323_6 ( .COUTX(na1323_3), .POUTX(na1323_6), .CINX(1'b0), .CINY1(na1322_4), .CINY2(na1322_5), .PINX(1'b0), .PINY1(na1322_7),
                      .PINY2(na1322_8), .OUT1(1'b0), .OUT2(na1323_2), .COMP_OUT(na1323_3_i) );
// C_AND///AND/      x35y45     80'h00_0078_12_0000_0C88_FFF0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1324_1 ( .OUT(na1324_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1324_4 ( .OUT(na1324_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1324_6 ( .COUTY1(na1324_4), .POUTY1(na1324_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1324_1), .OUT2(na1324_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x35y46     80'h00_0018_04_2056_5888_0CCF
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1325_1 ( .OUT(na1325_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(na1304_3), .CINY1(na1324_4), .PINX(1'b0), .PINY1(na1324_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1325_3 ( .COMP_OUT(na1325_3_i), .COMB1(na1325_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1325_6 ( .COUTY1(na1325_4), .COUTY2(na1325_5), .POUTY1(na1325_7), .CINX(na1304_3), .CINY1(na1324_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1324_7), .PINY2(1'b0), .OUT1(na1325_1), .OUT2(1'b0), .COMP_OUT(na1325_3_i) );
// C_MULTFa//O_O2//      x35y47     80'h00_0018_13_A477_34A6_0CCC
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1326_1 ( .COUTX(na1326_3), .COUTY1(na1326_4), .COUTY2(na1326_5), .POUTY1(na1326_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1305_3), .CINY1(na1325_4),
                      .CINY2(na1325_5), .PINX(1'b0), .PINY1(na1325_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x35y48     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1327_1 ( .OUT(na1327_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1326_4), .PINX(1'b0), .PINY1(na1326_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1327_3 ( .COMP_OUT(na1327_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1327_4 ( .OUT(na1327_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1326_4), .PINX(1'b0), .PINY1(na1326_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1327_6 ( .COUTX(na1327_3), .COUTY1(na1327_4), .COUTY2(na1327_5), .POUTY1(na1327_7), .POUTY2(na1327_8), .CINX(1'b0), .CINY1(na1326_4),
                      .CINY2(na1326_5), .PINX(1'b0), .PINY1(na1326_7), .PINY2(1'b0), .OUT1(na1327_1), .OUT2(na1327_2), .COMP_OUT(na1327_3_i) );
// C_MULT///MULT/      x35y49     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1328_1 ( .COUTY1(na1328_4), .COUTY2(na1328_5), .POUTY1(na1328_7), .POUTY2(na1328_8), .IN1(na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1307_3),
                      .CINY1(na1327_4), .CINY2(na1327_5), .PINX(na1307_6), .PINY1(na1327_7), .PINY2(na1327_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y50     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1329_1 ( .COUTX(na1329_3), .COUTY1(na1329_4), .COUTY2(na1329_5), .POUTX(na1329_6), .POUTY1(na1329_7), .POUTY2(na1329_8),
                      .IN1(~na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1308_3), .CINY1(na1328_4), .CINY2(na1328_5), .PINX(na1308_6), .PINY1(na1328_7), .PINY2(na1328_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y51     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1330_1 ( .COUTX(na1330_3), .COUTY1(na1330_4), .COUTY2(na1330_5), .POUTX(na1330_6), .POUTY1(na1330_7), .POUTY2(na1330_8),
                      .IN1(na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1309_3), .CINY1(na1329_4), .CINY2(na1329_5), .PINX(na1309_6), .PINY1(na1329_7), .PINY2(na1329_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y52     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1331_1 ( .COUTX(na1331_3), .COUTY1(na1331_4), .COUTY2(na1331_5), .POUTX(na1331_6), .POUTY1(na1331_7), .POUTY2(na1331_8),
                      .IN1(~na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1310_3), .CINY1(na1330_4), .CINY2(na1330_5), .PINX(na1310_6), .PINY1(na1330_7), .PINY2(na1330_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1332_1 ( .COUTX(na1332_3), .COUTY1(na1332_4), .COUTY2(na1332_5), .POUTX(na1332_6), .POUTY1(na1332_7), .POUTY2(na1332_8),
                      .IN1(na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1311_3), .CINY1(na1331_4), .CINY2(na1331_5), .PINX(na1311_6), .PINY1(na1331_7), .PINY2(na1331_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1333_1 ( .COUTX(na1333_3), .COUTY1(na1333_4), .COUTY2(na1333_5), .POUTX(na1333_6), .POUTY1(na1333_7), .POUTY2(na1333_8),
                      .IN1(~na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1312_3), .CINY1(na1332_4), .CINY2(na1332_5), .PINX(na1312_6), .PINY1(na1332_7), .PINY2(na1332_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1334_1 ( .COUTX(na1334_3), .COUTY1(na1334_4), .COUTY2(na1334_5), .POUTX(na1334_6), .POUTY1(na1334_7), .POUTY2(na1334_8),
                      .IN1(na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1313_3), .CINY1(na1333_4), .CINY2(na1333_5), .PINX(na1313_6), .PINY1(na1333_7), .PINY2(na1333_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1335_1 ( .COUTX(na1335_3), .COUTY1(na1335_4), .COUTY2(na1335_5), .POUTX(na1335_6), .POUTY1(na1335_7), .POUTY2(na1335_8),
                      .IN1(~na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1314_3), .CINY1(na1334_4), .CINY2(na1334_5), .PINX(na1314_6), .PINY1(na1334_7), .PINY2(na1334_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1336_1 ( .COUTX(na1336_3), .COUTY1(na1336_4), .COUTY2(na1336_5), .POUTX(na1336_6), .POUTY1(na1336_7), .POUTY2(na1336_8),
                      .IN1(na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1315_3), .CINY1(na1335_4), .CINY2(na1335_5), .PINX(na1315_6), .PINY1(na1335_7), .PINY2(na1335_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1337_1 ( .COUTX(na1337_3), .COUTY1(na1337_4), .COUTY2(na1337_5), .POUTX(na1337_6), .POUTY1(na1337_7), .POUTY2(na1337_8),
                      .IN1(~na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1316_3), .CINY1(na1336_4), .CINY2(na1336_5), .PINX(na1316_6), .PINY1(na1336_7), .PINY2(na1336_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1338_1 ( .COUTX(na1338_3), .COUTY1(na1338_4), .COUTY2(na1338_5), .POUTX(na1338_6), .POUTY1(na1338_7), .POUTY2(na1338_8),
                      .IN1(na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1317_3), .CINY1(na1337_4), .CINY2(na1337_5), .PINX(na1317_6), .PINY1(na1337_7), .PINY2(na1337_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1339_1 ( .COUTX(na1339_3), .COUTY1(na1339_4), .COUTY2(na1339_5), .POUTX(na1339_6), .POUTY1(na1339_7), .POUTY2(na1339_8),
                      .IN1(~na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1318_3), .CINY1(na1338_4), .CINY2(na1338_5), .PINX(na1318_6), .PINY1(na1338_7), .PINY2(na1338_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y61     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1340_1 ( .COUTX(na1340_3), .COUTY1(na1340_4), .COUTY2(na1340_5), .POUTX(na1340_6), .POUTY1(na1340_7), .POUTY2(na1340_8),
                      .IN1(na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1319_3), .CINY1(na1339_4), .CINY2(na1339_5), .PINX(na1319_6), .PINY1(na1339_7), .PINY2(na1339_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y62     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1341_1 ( .COUTX(na1341_3), .COUTY1(na1341_4), .COUTY2(na1341_5), .POUTX(na1341_6), .POUTY1(na1341_7), .POUTY2(na1341_8),
                      .IN1(~na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1320_3), .CINY1(na1340_4), .CINY2(na1340_5), .PINX(na1320_6), .PINY1(na1340_7), .PINY2(na1340_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y63     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1342_1 ( .COUTX(na1342_3), .COUTY1(na1342_4), .COUTY2(na1342_5), .POUTX(na1342_6), .POUTY1(na1342_7), .POUTY2(na1342_8),
                      .IN1(na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1321_3), .CINY1(na1341_4), .CINY2(na1341_5), .PINX(na1321_6), .PINY1(na1341_7), .PINY2(na1341_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y64     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1343_1 ( .COUTX(na1343_3), .COUTY1(na1343_4), .COUTY2(na1343_5), .POUTX(na1343_6), .POUTY1(na1343_7), .POUTY2(na1343_8),
                      .IN1(~na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1322_3), .CINY1(na1342_4), .CINY2(na1342_5), .PINX(na1322_6), .PINY1(na1342_7), .PINY2(na1342_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x35y65     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1344_1 ( .COUTX(na1344_3), .COUTY1(na1344_4), .COUTY2(na1344_5), .POUTX(na1344_6), .POUTY1(na1344_7), .POUTY2(na1344_8),
                      .IN1(na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1323_3), .CINY1(na1343_4), .CINY2(na1343_5), .PINX(na1323_6), .PINY1(na1343_7), .PINY2(na1343_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x35y66     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1345_3 ( .COMP_OUT(na1345_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1345_4 ( .OUT(na1345_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1344_4), .PINX(1'b0), .PINY1(na1344_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1345_6 ( .COUTX(na1345_3), .POUTX(na1345_6), .CINX(1'b0), .CINY1(na1344_4), .CINY2(na1344_5), .PINX(1'b0), .PINY1(na1344_7),
                      .PINY2(na1344_8), .OUT1(1'b0), .OUT2(na1345_2), .COMP_OUT(na1345_3_i) );
// C_AND///AND/      x36y46     80'h00_0078_12_0000_0C88_FFF0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1346_1 ( .OUT(na1346_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1346_4 ( .OUT(na1346_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1346_6 ( .COUTY1(na1346_4), .POUTY1(na1346_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1346_1), .OUT2(na1346_2), .COMP_OUT(1'b0) );
// C_OR//O_O1//      x36y47     80'h00_0018_04_2056_5EEE_0CC0
C_OR       #(.CPE_CFG (9'b0_0001_0110)) 
           _a1347_1 ( .OUT(na1347_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(na1326_3), .CINY1(na1346_4), .PINX(1'b0), .PINY1(na1346_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1347_3 ( .COMP_OUT(na1347_3_i), .COMB1(na1347_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1347_6 ( .COUTY1(na1347_4), .COUTY2(na1347_5), .POUTY1(na1347_7), .CINX(na1326_3), .CINY1(na1346_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1346_7), .PINY2(1'b0), .OUT1(na1347_1), .OUT2(1'b0), .COMP_OUT(na1347_3_i) );
// C_MULTFb//O_O2//      x36y48     80'h00_0018_13_A477_3EA6_0CCC
C_MULTFb   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1348_1 ( .COUTX(na1348_3), .COUTY1(na1348_4), .COUTY2(na1348_5), .POUTY1(na1348_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1327_3), .CINY1(na1347_4),
                      .CINY2(na1347_5), .PINX(1'b0), .PINY1(na1347_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_O2/AND/      x36y49     80'h00_0078_35_A471_3C88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1349_1 ( .OUT(na1349_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1348_4), .PINX(1'b0), .PINY1(na1348_7) );
C_O_O2     #(.CPE_CFG ()) 
           _a1349_3 ( .COMP_OUT(na1349_3_i), .COMB1(1'b0), .COMB2(na1349_2) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1349_4 ( .OUT(na1349_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1348_4), .PINX(1'b0), .PINY1(na1348_7) );
C_CPlines  #(.CPE_CFG (19'h3_5A47)) 
           _a1349_6 ( .COUTX(na1349_3), .COUTY1(na1349_4), .COUTY2(na1349_5), .POUTY1(na1349_7), .POUTY2(na1349_8), .CINX(1'b0), .CINY1(na1348_4),
                      .CINY2(na1348_5), .PINX(1'b0), .PINY1(na1348_7), .PINY2(1'b0), .OUT1(na1349_1), .OUT2(na1349_2), .COMP_OUT(na1349_3_i) );
// C_MULT///MULT/      x36y50     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1350_1 ( .COUTY1(na1350_4), .COUTY2(na1350_5), .POUTY1(na1350_7), .POUTY2(na1350_8), .IN1(~na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1329_3),
                      .CINY1(na1349_4), .CINY2(na1349_5), .PINX(na1329_6), .PINY1(na1349_7), .PINY2(na1349_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y51     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1351_1 ( .COUTX(na1351_3), .COUTY1(na1351_4), .COUTY2(na1351_5), .POUTX(na1351_6), .POUTY1(na1351_7), .POUTY2(na1351_8),
                      .IN1(na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1330_3), .CINY1(na1350_4), .CINY2(na1350_5), .PINX(na1330_6), .PINY1(na1350_7), .PINY2(na1350_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y52     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1352_1 ( .COUTX(na1352_3), .COUTY1(na1352_4), .COUTY2(na1352_5), .POUTX(na1352_6), .POUTY1(na1352_7), .POUTY2(na1352_8),
                      .IN1(~na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1331_3), .CINY1(na1351_4), .CINY2(na1351_5), .PINX(na1331_6), .PINY1(na1351_7), .PINY2(na1351_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1353_1 ( .COUTX(na1353_3), .COUTY1(na1353_4), .COUTY2(na1353_5), .POUTX(na1353_6), .POUTY1(na1353_7), .POUTY2(na1353_8),
                      .IN1(na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1332_3), .CINY1(na1352_4), .CINY2(na1352_5), .PINX(na1332_6), .PINY1(na1352_7), .PINY2(na1352_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1354_1 ( .COUTX(na1354_3), .COUTY1(na1354_4), .COUTY2(na1354_5), .POUTX(na1354_6), .POUTY1(na1354_7), .POUTY2(na1354_8),
                      .IN1(~na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1333_3), .CINY1(na1353_4), .CINY2(na1353_5), .PINX(na1333_6), .PINY1(na1353_7), .PINY2(na1353_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1355_1 ( .COUTX(na1355_3), .COUTY1(na1355_4), .COUTY2(na1355_5), .POUTX(na1355_6), .POUTY1(na1355_7), .POUTY2(na1355_8),
                      .IN1(na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1334_3), .CINY1(na1354_4), .CINY2(na1354_5), .PINX(na1334_6), .PINY1(na1354_7), .PINY2(na1354_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1356_1 ( .COUTX(na1356_3), .COUTY1(na1356_4), .COUTY2(na1356_5), .POUTX(na1356_6), .POUTY1(na1356_7), .POUTY2(na1356_8),
                      .IN1(~na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1335_3), .CINY1(na1355_4), .CINY2(na1355_5), .PINX(na1335_6), .PINY1(na1355_7), .PINY2(na1355_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1357_1 ( .COUTX(na1357_3), .COUTY1(na1357_4), .COUTY2(na1357_5), .POUTX(na1357_6), .POUTY1(na1357_7), .POUTY2(na1357_8),
                      .IN1(na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1336_3), .CINY1(na1356_4), .CINY2(na1356_5), .PINX(na1336_6), .PINY1(na1356_7), .PINY2(na1356_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1358_1 ( .COUTX(na1358_3), .COUTY1(na1358_4), .COUTY2(na1358_5), .POUTX(na1358_6), .POUTY1(na1358_7), .POUTY2(na1358_8),
                      .IN1(~na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1337_3), .CINY1(na1357_4), .CINY2(na1357_5), .PINX(na1337_6), .PINY1(na1357_7), .PINY2(na1357_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1359_1 ( .COUTX(na1359_3), .COUTY1(na1359_4), .COUTY2(na1359_5), .POUTX(na1359_6), .POUTY1(na1359_7), .POUTY2(na1359_8),
                      .IN1(na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1338_3), .CINY1(na1358_4), .CINY2(na1358_5), .PINX(na1338_6), .PINY1(na1358_7), .PINY2(na1358_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1360_1 ( .COUTX(na1360_3), .COUTY1(na1360_4), .COUTY2(na1360_5), .POUTX(na1360_6), .POUTY1(na1360_7), .POUTY2(na1360_8),
                      .IN1(~na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1339_3), .CINY1(na1359_4), .CINY2(na1359_5), .PINX(na1339_6), .PINY1(na1359_7), .PINY2(na1359_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y61     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1361_1 ( .COUTX(na1361_3), .COUTY1(na1361_4), .COUTY2(na1361_5), .POUTX(na1361_6), .POUTY1(na1361_7), .POUTY2(na1361_8),
                      .IN1(na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1340_3), .CINY1(na1360_4), .CINY2(na1360_5), .PINX(na1340_6), .PINY1(na1360_7), .PINY2(na1360_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y62     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1362_1 ( .COUTX(na1362_3), .COUTY1(na1362_4), .COUTY2(na1362_5), .POUTX(na1362_6), .POUTY1(na1362_7), .POUTY2(na1362_8),
                      .IN1(~na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1341_3), .CINY1(na1361_4), .CINY2(na1361_5), .PINX(na1341_6), .PINY1(na1361_7), .PINY2(na1361_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y63     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1363_1 ( .COUTX(na1363_3), .COUTY1(na1363_4), .COUTY2(na1363_5), .POUTX(na1363_6), .POUTY1(na1363_7), .POUTY2(na1363_8),
                      .IN1(na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1342_3), .CINY1(na1362_4), .CINY2(na1362_5), .PINX(na1342_6), .PINY1(na1362_7), .PINY2(na1362_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y64     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1364_1 ( .COUTX(na1364_3), .COUTY1(na1364_4), .COUTY2(na1364_5), .POUTX(na1364_6), .POUTY1(na1364_7), .POUTY2(na1364_8),
                      .IN1(~na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1343_3), .CINY1(na1363_4), .CINY2(na1363_5), .PINX(na1343_6), .PINY1(na1363_7), .PINY2(na1363_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y65     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1365_1 ( .COUTX(na1365_3), .COUTY1(na1365_4), .COUTY2(na1365_5), .POUTX(na1365_6), .POUTY1(na1365_7), .POUTY2(na1365_8),
                      .IN1(na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1344_3), .CINY1(na1364_4), .CINY2(na1364_5), .PINX(na1344_6), .PINY1(na1364_7), .PINY2(na1364_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x36y66     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1366_1 ( .COUTX(na1366_3), .COUTY1(na1366_4), .COUTY2(na1366_5), .POUTX(na1366_6), .POUTY1(na1366_7), .POUTY2(na1366_8),
                      .IN1(~na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1345_3), .CINY1(na1365_4), .CINY2(na1365_5), .PINX(na1345_6), .PINY1(na1365_7), .PINY2(na1365_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x36y67     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1367_3 ( .COMP_OUT(na1367_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1367_4 ( .OUT(na1367_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1366_4), .PINX(1'b0), .PINY1(na1366_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1367_6 ( .COUTX(na1367_3), .POUTX(na1367_6), .CINX(1'b0), .CINY1(na1366_4), .CINY2(na1366_5), .PINX(1'b0), .PINY1(na1366_7),
                      .PINY2(na1366_8), .OUT1(1'b0), .OUT2(na1367_2), .COMP_OUT(na1367_3_i) );
// C_AND///AND/      x37y47     80'h00_0078_12_0000_0C88_FFF0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1368_1 ( .OUT(na1368_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1368_4 ( .OUT(na1368_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1368_6 ( .COUTY1(na1368_4), .POUTY1(na1368_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1368_1), .OUT2(na1368_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x37y48     80'h00_0018_04_2056_5888_0CCF
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1369_1 ( .OUT(na1369_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(na1348_3), .CINY1(na1368_4), .PINX(1'b0), .PINY1(na1368_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1369_3 ( .COMP_OUT(na1369_3_i), .COMB1(na1369_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1369_6 ( .COUTY1(na1369_4), .COUTY2(na1369_5), .POUTY1(na1369_7), .CINX(na1348_3), .CINY1(na1368_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1368_7), .PINY2(1'b0), .OUT1(na1369_1), .OUT2(1'b0), .COMP_OUT(na1369_3_i) );
// C_MULTFa//O_O2//      x37y49     80'h00_0018_13_A477_34A6_0CCC
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1370_1 ( .COUTX(na1370_3), .COUTY1(na1370_4), .COUTY2(na1370_5), .POUTY1(na1370_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1349_3), .CINY1(na1369_4),
                      .CINY2(na1369_5), .PINX(1'b0), .PINY1(na1369_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x37y50     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1371_1 ( .OUT(na1371_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1370_4), .PINX(1'b0), .PINY1(na1370_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1371_3 ( .COMP_OUT(na1371_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1371_4 ( .OUT(na1371_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1370_4), .PINX(1'b0), .PINY1(na1370_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1371_6 ( .COUTX(na1371_3), .COUTY1(na1371_4), .COUTY2(na1371_5), .POUTY1(na1371_7), .POUTY2(na1371_8), .CINX(1'b0), .CINY1(na1370_4),
                      .CINY2(na1370_5), .PINX(1'b0), .PINY1(na1370_7), .PINY2(1'b0), .OUT1(na1371_1), .OUT2(na1371_2), .COMP_OUT(na1371_3_i) );
// C_MULT///MULT/      x37y51     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1372_1 ( .COUTY1(na1372_4), .COUTY2(na1372_5), .POUTY1(na1372_7), .POUTY2(na1372_8), .IN1(na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1351_3),
                      .CINY1(na1371_4), .CINY2(na1371_5), .PINX(na1351_6), .PINY1(na1371_7), .PINY2(na1371_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y52     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1373_1 ( .COUTX(na1373_3), .COUTY1(na1373_4), .COUTY2(na1373_5), .POUTX(na1373_6), .POUTY1(na1373_7), .POUTY2(na1373_8),
                      .IN1(~na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1352_3), .CINY1(na1372_4), .CINY2(na1372_5), .PINX(na1352_6), .PINY1(na1372_7), .PINY2(na1372_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1374_1 ( .COUTX(na1374_3), .COUTY1(na1374_4), .COUTY2(na1374_5), .POUTX(na1374_6), .POUTY1(na1374_7), .POUTY2(na1374_8),
                      .IN1(na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1353_3), .CINY1(na1373_4), .CINY2(na1373_5), .PINX(na1353_6), .PINY1(na1373_7), .PINY2(na1373_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1375_1 ( .COUTX(na1375_3), .COUTY1(na1375_4), .COUTY2(na1375_5), .POUTX(na1375_6), .POUTY1(na1375_7), .POUTY2(na1375_8),
                      .IN1(~na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1354_3), .CINY1(na1374_4), .CINY2(na1374_5), .PINX(na1354_6), .PINY1(na1374_7), .PINY2(na1374_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1376_1 ( .COUTX(na1376_3), .COUTY1(na1376_4), .COUTY2(na1376_5), .POUTX(na1376_6), .POUTY1(na1376_7), .POUTY2(na1376_8),
                      .IN1(na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1355_3), .CINY1(na1375_4), .CINY2(na1375_5), .PINX(na1355_6), .PINY1(na1375_7), .PINY2(na1375_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1377_1 ( .COUTX(na1377_3), .COUTY1(na1377_4), .COUTY2(na1377_5), .POUTX(na1377_6), .POUTY1(na1377_7), .POUTY2(na1377_8),
                      .IN1(~na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1356_3), .CINY1(na1376_4), .CINY2(na1376_5), .PINX(na1356_6), .PINY1(na1376_7), .PINY2(na1376_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1378_1 ( .COUTX(na1378_3), .COUTY1(na1378_4), .COUTY2(na1378_5), .POUTX(na1378_6), .POUTY1(na1378_7), .POUTY2(na1378_8),
                      .IN1(na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1357_3), .CINY1(na1377_4), .CINY2(na1377_5), .PINX(na1357_6), .PINY1(na1377_7), .PINY2(na1377_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1379_1 ( .COUTX(na1379_3), .COUTY1(na1379_4), .COUTY2(na1379_5), .POUTX(na1379_6), .POUTY1(na1379_7), .POUTY2(na1379_8),
                      .IN1(~na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1358_3), .CINY1(na1378_4), .CINY2(na1378_5), .PINX(na1358_6), .PINY1(na1378_7), .PINY2(na1378_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1380_1 ( .COUTX(na1380_3), .COUTY1(na1380_4), .COUTY2(na1380_5), .POUTX(na1380_6), .POUTY1(na1380_7), .POUTY2(na1380_8),
                      .IN1(na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1359_3), .CINY1(na1379_4), .CINY2(na1379_5), .PINX(na1359_6), .PINY1(na1379_7), .PINY2(na1379_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1381_1 ( .COUTX(na1381_3), .COUTY1(na1381_4), .COUTY2(na1381_5), .POUTX(na1381_6), .POUTY1(na1381_7), .POUTY2(na1381_8),
                      .IN1(~na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1360_3), .CINY1(na1380_4), .CINY2(na1380_5), .PINX(na1360_6), .PINY1(na1380_7), .PINY2(na1380_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y61     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1382_1 ( .COUTX(na1382_3), .COUTY1(na1382_4), .COUTY2(na1382_5), .POUTX(na1382_6), .POUTY1(na1382_7), .POUTY2(na1382_8),
                      .IN1(na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1361_3), .CINY1(na1381_4), .CINY2(na1381_5), .PINX(na1361_6), .PINY1(na1381_7), .PINY2(na1381_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y62     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1383_1 ( .COUTX(na1383_3), .COUTY1(na1383_4), .COUTY2(na1383_5), .POUTX(na1383_6), .POUTY1(na1383_7), .POUTY2(na1383_8),
                      .IN1(~na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1362_3), .CINY1(na1382_4), .CINY2(na1382_5), .PINX(na1362_6), .PINY1(na1382_7), .PINY2(na1382_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y63     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1384_1 ( .COUTX(na1384_3), .COUTY1(na1384_4), .COUTY2(na1384_5), .POUTX(na1384_6), .POUTY1(na1384_7), .POUTY2(na1384_8),
                      .IN1(na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1363_3), .CINY1(na1383_4), .CINY2(na1383_5), .PINX(na1363_6), .PINY1(na1383_7), .PINY2(na1383_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y64     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1385_1 ( .COUTX(na1385_3), .COUTY1(na1385_4), .COUTY2(na1385_5), .POUTX(na1385_6), .POUTY1(na1385_7), .POUTY2(na1385_8),
                      .IN1(~na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1364_3), .CINY1(na1384_4), .CINY2(na1384_5), .PINX(na1364_6), .PINY1(na1384_7), .PINY2(na1384_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y65     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1386_1 ( .COUTX(na1386_3), .COUTY1(na1386_4), .COUTY2(na1386_5), .POUTX(na1386_6), .POUTY1(na1386_7), .POUTY2(na1386_8),
                      .IN1(na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1365_3), .CINY1(na1385_4), .CINY2(na1385_5), .PINX(na1365_6), .PINY1(na1385_7), .PINY2(na1385_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y66     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1387_1 ( .COUTX(na1387_3), .COUTY1(na1387_4), .COUTY2(na1387_5), .POUTX(na1387_6), .POUTY1(na1387_7), .POUTY2(na1387_8),
                      .IN1(~na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1366_3), .CINY1(na1386_4), .CINY2(na1386_5), .PINX(na1366_6), .PINY1(na1386_7), .PINY2(na1386_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x37y67     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1388_1 ( .COUTX(na1388_3), .COUTY1(na1388_4), .COUTY2(na1388_5), .POUTX(na1388_6), .POUTY1(na1388_7), .POUTY2(na1388_8),
                      .IN1(na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1367_3), .CINY1(na1387_4), .CINY2(na1387_5), .PINX(na1367_6), .PINY1(na1387_7), .PINY2(na1387_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x37y68     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1389_3 ( .COMP_OUT(na1389_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1389_4 ( .OUT(na1389_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1388_4), .PINX(1'b0), .PINY1(na1388_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1389_6 ( .COUTX(na1389_3), .POUTX(na1389_6), .CINX(1'b0), .CINY1(na1388_4), .CINY2(na1388_5), .PINX(1'b0), .PINY1(na1388_7),
                      .PINY2(na1388_8), .OUT1(1'b0), .OUT2(na1389_2), .COMP_OUT(na1389_3_i) );
// C_AND///AND/      x38y48     80'h00_0078_12_0000_0C88_F0FF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1390_1 ( .OUT(na1390_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1390_4 ( .OUT(na1390_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1390_6 ( .COUTY1(na1390_4), .POUTY1(na1390_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1390_1), .OUT2(na1390_2), .COMP_OUT(1'b0) );
// C_OR//O_O1//      x38y49     80'h00_0018_04_2056_5EEE_0CC0
C_OR       #(.CPE_CFG (9'b0_0001_0110)) 
           _a1391_1 ( .OUT(na1391_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(na1370_3), .CINY1(na1390_4), .PINX(1'b0), .PINY1(na1390_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1391_3 ( .COMP_OUT(na1391_3_i), .COMB1(na1391_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1391_6 ( .COUTY1(na1391_4), .COUTY2(na1391_5), .POUTY1(na1391_7), .CINX(na1370_3), .CINY1(na1390_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1390_7), .PINY2(1'b0), .OUT1(na1391_1), .OUT2(1'b0), .COMP_OUT(na1391_3_i) );
// C_MULTFb//O_O2//      x38y50     80'h00_0018_13_A477_3EA6_0CCC
C_MULTFb   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1392_1 ( .COUTX(na1392_3), .COUTY1(na1392_4), .COUTY2(na1392_5), .POUTY1(na1392_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1371_3), .CINY1(na1391_4),
                      .CINY2(na1391_5), .PINX(1'b0), .PINY1(na1391_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_O2/AND/      x38y51     80'h00_0078_35_A471_3C88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1393_1 ( .OUT(na1393_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1392_4), .PINX(1'b0), .PINY1(na1392_7) );
C_O_O2     #(.CPE_CFG ()) 
           _a1393_3 ( .COMP_OUT(na1393_3_i), .COMB1(1'b0), .COMB2(na1393_2) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1393_4 ( .OUT(na1393_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1392_4), .PINX(1'b0), .PINY1(na1392_7) );
C_CPlines  #(.CPE_CFG (19'h3_5A47)) 
           _a1393_6 ( .COUTX(na1393_3), .COUTY1(na1393_4), .COUTY2(na1393_5), .POUTY1(na1393_7), .POUTY2(na1393_8), .CINX(1'b0), .CINY1(na1392_4),
                      .CINY2(na1392_5), .PINX(1'b0), .PINY1(na1392_7), .PINY2(1'b0), .OUT1(na1393_1), .OUT2(na1393_2), .COMP_OUT(na1393_3_i) );
// C_MULT///MULT/      x38y52     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1394_1 ( .COUTY1(na1394_4), .COUTY2(na1394_5), .POUTY1(na1394_7), .POUTY2(na1394_8), .IN1(~na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1373_3),
                      .CINY1(na1393_4), .CINY2(na1393_5), .PINX(na1373_6), .PINY1(na1393_7), .PINY2(na1393_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y53     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1395_1 ( .COUTX(na1395_3), .COUTY1(na1395_4), .COUTY2(na1395_5), .POUTX(na1395_6), .POUTY1(na1395_7), .POUTY2(na1395_8),
                      .IN1(na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1374_3), .CINY1(na1394_4), .CINY2(na1394_5), .PINX(na1374_6), .PINY1(na1394_7), .PINY2(na1394_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1396_1 ( .COUTX(na1396_3), .COUTY1(na1396_4), .COUTY2(na1396_5), .POUTX(na1396_6), .POUTY1(na1396_7), .POUTY2(na1396_8),
                      .IN1(~na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1375_3), .CINY1(na1395_4), .CINY2(na1395_5), .PINX(na1375_6), .PINY1(na1395_7), .PINY2(na1395_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1397_1 ( .COUTX(na1397_3), .COUTY1(na1397_4), .COUTY2(na1397_5), .POUTX(na1397_6), .POUTY1(na1397_7), .POUTY2(na1397_8),
                      .IN1(na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1376_3), .CINY1(na1396_4), .CINY2(na1396_5), .PINX(na1376_6), .PINY1(na1396_7), .PINY2(na1396_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1398_1 ( .COUTX(na1398_3), .COUTY1(na1398_4), .COUTY2(na1398_5), .POUTX(na1398_6), .POUTY1(na1398_7), .POUTY2(na1398_8),
                      .IN1(~na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1377_3), .CINY1(na1397_4), .CINY2(na1397_5), .PINX(na1377_6), .PINY1(na1397_7), .PINY2(na1397_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1399_1 ( .COUTX(na1399_3), .COUTY1(na1399_4), .COUTY2(na1399_5), .POUTX(na1399_6), .POUTY1(na1399_7), .POUTY2(na1399_8),
                      .IN1(na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1378_3), .CINY1(na1398_4), .CINY2(na1398_5), .PINX(na1378_6), .PINY1(na1398_7), .PINY2(na1398_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1400_1 ( .COUTX(na1400_3), .COUTY1(na1400_4), .COUTY2(na1400_5), .POUTX(na1400_6), .POUTY1(na1400_7), .POUTY2(na1400_8),
                      .IN1(~na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1379_3), .CINY1(na1399_4), .CINY2(na1399_5), .PINX(na1379_6), .PINY1(na1399_7), .PINY2(na1399_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1401_1 ( .COUTX(na1401_3), .COUTY1(na1401_4), .COUTY2(na1401_5), .POUTX(na1401_6), .POUTY1(na1401_7), .POUTY2(na1401_8),
                      .IN1(na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1380_3), .CINY1(na1400_4), .CINY2(na1400_5), .PINX(na1380_6), .PINY1(na1400_7), .PINY2(na1400_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1402_1 ( .COUTX(na1402_3), .COUTY1(na1402_4), .COUTY2(na1402_5), .POUTX(na1402_6), .POUTY1(na1402_7), .POUTY2(na1402_8),
                      .IN1(~na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1381_3), .CINY1(na1401_4), .CINY2(na1401_5), .PINX(na1381_6), .PINY1(na1401_7), .PINY2(na1401_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y61     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1403_1 ( .COUTX(na1403_3), .COUTY1(na1403_4), .COUTY2(na1403_5), .POUTX(na1403_6), .POUTY1(na1403_7), .POUTY2(na1403_8),
                      .IN1(na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1382_3), .CINY1(na1402_4), .CINY2(na1402_5), .PINX(na1382_6), .PINY1(na1402_7), .PINY2(na1402_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y62     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1404_1 ( .COUTX(na1404_3), .COUTY1(na1404_4), .COUTY2(na1404_5), .POUTX(na1404_6), .POUTY1(na1404_7), .POUTY2(na1404_8),
                      .IN1(~na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1383_3), .CINY1(na1403_4), .CINY2(na1403_5), .PINX(na1383_6), .PINY1(na1403_7), .PINY2(na1403_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y63     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1405_1 ( .COUTX(na1405_3), .COUTY1(na1405_4), .COUTY2(na1405_5), .POUTX(na1405_6), .POUTY1(na1405_7), .POUTY2(na1405_8),
                      .IN1(na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1384_3), .CINY1(na1404_4), .CINY2(na1404_5), .PINX(na1384_6), .PINY1(na1404_7), .PINY2(na1404_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y64     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1406_1 ( .COUTX(na1406_3), .COUTY1(na1406_4), .COUTY2(na1406_5), .POUTX(na1406_6), .POUTY1(na1406_7), .POUTY2(na1406_8),
                      .IN1(~na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1385_3), .CINY1(na1405_4), .CINY2(na1405_5), .PINX(na1385_6), .PINY1(na1405_7), .PINY2(na1405_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y65     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1407_1 ( .COUTX(na1407_3), .COUTY1(na1407_4), .COUTY2(na1407_5), .POUTX(na1407_6), .POUTY1(na1407_7), .POUTY2(na1407_8),
                      .IN1(na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1386_3), .CINY1(na1406_4), .CINY2(na1406_5), .PINX(na1386_6), .PINY1(na1406_7), .PINY2(na1406_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y66     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1408_1 ( .COUTX(na1408_3), .COUTY1(na1408_4), .COUTY2(na1408_5), .POUTX(na1408_6), .POUTY1(na1408_7), .POUTY2(na1408_8),
                      .IN1(~na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1387_3), .CINY1(na1407_4), .CINY2(na1407_5), .PINX(na1387_6), .PINY1(na1407_7), .PINY2(na1407_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y67     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1409_1 ( .COUTX(na1409_3), .COUTY1(na1409_4), .COUTY2(na1409_5), .POUTX(na1409_6), .POUTY1(na1409_7), .POUTY2(na1409_8),
                      .IN1(na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1388_3), .CINY1(na1408_4), .CINY2(na1408_5), .PINX(na1388_6), .PINY1(na1408_7), .PINY2(na1408_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x38y68     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1410_1 ( .COUTX(na1410_3), .COUTY1(na1410_4), .COUTY2(na1410_5), .POUTX(na1410_6), .POUTY1(na1410_7), .POUTY2(na1410_8),
                      .IN1(~na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1389_3), .CINY1(na1409_4), .CINY2(na1409_5), .PINX(na1389_6), .PINY1(na1409_7), .PINY2(na1409_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x38y69     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1411_3 ( .COMP_OUT(na1411_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1411_4 ( .OUT(na1411_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1410_4), .PINX(1'b0), .PINY1(na1410_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1411_6 ( .COUTX(na1411_3), .POUTX(na1411_6), .CINX(1'b0), .CINY1(na1410_4), .CINY2(na1410_5), .PINX(1'b0), .PINY1(na1410_7),
                      .PINY2(na1410_8), .OUT1(1'b0), .OUT2(na1411_2), .COMP_OUT(na1411_3_i) );
// C_AND///AND/      x39y49     80'h00_0078_12_0000_0C88_FFFF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1412_1 ( .OUT(na1412_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1412_4 ( .OUT(na1412_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1412_6 ( .COUTY1(na1412_4), .POUTY1(na1412_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1412_1), .OUT2(na1412_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x39y50     80'h00_0018_04_2056_5888_0CCF
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1413_1 ( .OUT(na1413_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(na1392_3), .CINY1(na1412_4), .PINX(1'b0), .PINY1(na1412_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1413_3 ( .COMP_OUT(na1413_3_i), .COMB1(na1413_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1413_6 ( .COUTY1(na1413_4), .COUTY2(na1413_5), .POUTY1(na1413_7), .CINX(na1392_3), .CINY1(na1412_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1412_7), .PINY2(1'b0), .OUT1(na1413_1), .OUT2(1'b0), .COMP_OUT(na1413_3_i) );
// C_MULTFa//O_O2//      x39y51     80'h00_0018_13_A477_34A6_0CCC
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1414_1 ( .COUTX(na1414_3), .COUTY1(na1414_4), .COUTY2(na1414_5), .POUTY1(na1414_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1393_3), .CINY1(na1413_4),
                      .CINY2(na1413_5), .PINX(1'b0), .PINY1(na1413_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x39y52     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1415_1 ( .OUT(na1415_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1414_4), .PINX(1'b0), .PINY1(na1414_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1415_3 ( .COMP_OUT(na1415_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1415_4 ( .OUT(na1415_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1414_4), .PINX(1'b0), .PINY1(na1414_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1415_6 ( .COUTX(na1415_3), .COUTY1(na1415_4), .COUTY2(na1415_5), .POUTY1(na1415_7), .POUTY2(na1415_8), .CINX(1'b0), .CINY1(na1414_4),
                      .CINY2(na1414_5), .PINX(1'b0), .PINY1(na1414_7), .PINY2(1'b0), .OUT1(na1415_1), .OUT2(na1415_2), .COMP_OUT(na1415_3_i) );
// C_MULT///MULT/      x39y53     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1416_1 ( .COUTY1(na1416_4), .COUTY2(na1416_5), .POUTY1(na1416_7), .POUTY2(na1416_8), .IN1(na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1395_3),
                      .CINY1(na1415_4), .CINY2(na1415_5), .PINX(na1395_6), .PINY1(na1415_7), .PINY2(na1415_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y54     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1417_1 ( .COUTX(na1417_3), .COUTY1(na1417_4), .COUTY2(na1417_5), .POUTX(na1417_6), .POUTY1(na1417_7), .POUTY2(na1417_8),
                      .IN1(~na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1396_3), .CINY1(na1416_4), .CINY2(na1416_5), .PINX(na1396_6), .PINY1(na1416_7), .PINY2(na1416_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1418_1 ( .COUTX(na1418_3), .COUTY1(na1418_4), .COUTY2(na1418_5), .POUTX(na1418_6), .POUTY1(na1418_7), .POUTY2(na1418_8),
                      .IN1(na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1397_3), .CINY1(na1417_4), .CINY2(na1417_5), .PINX(na1397_6), .PINY1(na1417_7), .PINY2(na1417_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1419_1 ( .COUTX(na1419_3), .COUTY1(na1419_4), .COUTY2(na1419_5), .POUTX(na1419_6), .POUTY1(na1419_7), .POUTY2(na1419_8),
                      .IN1(~na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1398_3), .CINY1(na1418_4), .CINY2(na1418_5), .PINX(na1398_6), .PINY1(na1418_7), .PINY2(na1418_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1420_1 ( .COUTX(na1420_3), .COUTY1(na1420_4), .COUTY2(na1420_5), .POUTX(na1420_6), .POUTY1(na1420_7), .POUTY2(na1420_8),
                      .IN1(na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1399_3), .CINY1(na1419_4), .CINY2(na1419_5), .PINX(na1399_6), .PINY1(na1419_7), .PINY2(na1419_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1421_1 ( .COUTX(na1421_3), .COUTY1(na1421_4), .COUTY2(na1421_5), .POUTX(na1421_6), .POUTY1(na1421_7), .POUTY2(na1421_8),
                      .IN1(~na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1400_3), .CINY1(na1420_4), .CINY2(na1420_5), .PINX(na1400_6), .PINY1(na1420_7), .PINY2(na1420_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1422_1 ( .COUTX(na1422_3), .COUTY1(na1422_4), .COUTY2(na1422_5), .POUTX(na1422_6), .POUTY1(na1422_7), .POUTY2(na1422_8),
                      .IN1(na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1401_3), .CINY1(na1421_4), .CINY2(na1421_5), .PINX(na1401_6), .PINY1(na1421_7), .PINY2(na1421_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1423_1 ( .COUTX(na1423_3), .COUTY1(na1423_4), .COUTY2(na1423_5), .POUTX(na1423_6), .POUTY1(na1423_7), .POUTY2(na1423_8),
                      .IN1(~na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1402_3), .CINY1(na1422_4), .CINY2(na1422_5), .PINX(na1402_6), .PINY1(na1422_7), .PINY2(na1422_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y61     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1424_1 ( .COUTX(na1424_3), .COUTY1(na1424_4), .COUTY2(na1424_5), .POUTX(na1424_6), .POUTY1(na1424_7), .POUTY2(na1424_8),
                      .IN1(na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1403_3), .CINY1(na1423_4), .CINY2(na1423_5), .PINX(na1403_6), .PINY1(na1423_7), .PINY2(na1423_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y62     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1425_1 ( .COUTX(na1425_3), .COUTY1(na1425_4), .COUTY2(na1425_5), .POUTX(na1425_6), .POUTY1(na1425_7), .POUTY2(na1425_8),
                      .IN1(~na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1404_3), .CINY1(na1424_4), .CINY2(na1424_5), .PINX(na1404_6), .PINY1(na1424_7), .PINY2(na1424_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y63     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1426_1 ( .COUTX(na1426_3), .COUTY1(na1426_4), .COUTY2(na1426_5), .POUTX(na1426_6), .POUTY1(na1426_7), .POUTY2(na1426_8),
                      .IN1(na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1405_3), .CINY1(na1425_4), .CINY2(na1425_5), .PINX(na1405_6), .PINY1(na1425_7), .PINY2(na1425_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y64     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1427_1 ( .COUTX(na1427_3), .COUTY1(na1427_4), .COUTY2(na1427_5), .POUTX(na1427_6), .POUTY1(na1427_7), .POUTY2(na1427_8),
                      .IN1(~na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1406_3), .CINY1(na1426_4), .CINY2(na1426_5), .PINX(na1406_6), .PINY1(na1426_7), .PINY2(na1426_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y65     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1428_1 ( .COUTX(na1428_3), .COUTY1(na1428_4), .COUTY2(na1428_5), .POUTX(na1428_6), .POUTY1(na1428_7), .POUTY2(na1428_8),
                      .IN1(na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1407_3), .CINY1(na1427_4), .CINY2(na1427_5), .PINX(na1407_6), .PINY1(na1427_7), .PINY2(na1427_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y66     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1429_1 ( .COUTX(na1429_3), .COUTY1(na1429_4), .COUTY2(na1429_5), .POUTX(na1429_6), .POUTY1(na1429_7), .POUTY2(na1429_8),
                      .IN1(~na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1408_3), .CINY1(na1428_4), .CINY2(na1428_5), .PINX(na1408_6), .PINY1(na1428_7), .PINY2(na1428_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y67     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1430_1 ( .COUTX(na1430_3), .COUTY1(na1430_4), .COUTY2(na1430_5), .POUTX(na1430_6), .POUTY1(na1430_7), .POUTY2(na1430_8),
                      .IN1(na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1409_3), .CINY1(na1429_4), .CINY2(na1429_5), .PINX(na1409_6), .PINY1(na1429_7), .PINY2(na1429_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y68     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1431_1 ( .COUTX(na1431_3), .COUTY1(na1431_4), .COUTY2(na1431_5), .POUTX(na1431_6), .POUTY1(na1431_7), .POUTY2(na1431_8),
                      .IN1(~na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1410_3), .CINY1(na1430_4), .CINY2(na1430_5), .PINX(na1410_6), .PINY1(na1430_7), .PINY2(na1430_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x39y69     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1432_1 ( .COUTX(na1432_3), .COUTY1(na1432_4), .COUTY2(na1432_5), .POUTX(na1432_6), .POUTY1(na1432_7), .POUTY2(na1432_8),
                      .IN1(na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1411_3), .CINY1(na1431_4), .CINY2(na1431_5), .PINX(na1411_6), .PINY1(na1431_7), .PINY2(na1431_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x39y70     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1433_3 ( .COMP_OUT(na1433_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1433_4 ( .OUT(na1433_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1432_4), .PINX(1'b0), .PINY1(na1432_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1433_6 ( .COUTX(na1433_3), .POUTX(na1433_6), .CINX(1'b0), .CINY1(na1432_4), .CINY2(na1432_5), .PINX(1'b0), .PINY1(na1432_7),
                      .PINY2(na1432_8), .OUT1(1'b0), .OUT2(na1433_2), .COMP_OUT(na1433_3_i) );
// C_AND///AND/      x40y50     80'h00_0078_12_0000_0C88_FFF0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1434_1 ( .OUT(na1434_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1434_4 ( .OUT(na1434_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1434_6 ( .COUTY1(na1434_4), .POUTY1(na1434_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1434_1), .OUT2(na1434_2), .COMP_OUT(1'b0) );
// C_OR//O_O1//      x40y51     80'h00_0018_04_2056_5EEE_0CC0
C_OR       #(.CPE_CFG (9'b0_0001_0110)) 
           _a1435_1 ( .OUT(na1435_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(na1414_3), .CINY1(na1434_4), .PINX(1'b0), .PINY1(na1434_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1435_3 ( .COMP_OUT(na1435_3_i), .COMB1(na1435_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1435_6 ( .COUTY1(na1435_4), .COUTY2(na1435_5), .POUTY1(na1435_7), .CINX(na1414_3), .CINY1(na1434_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1434_7), .PINY2(1'b0), .OUT1(na1435_1), .OUT2(1'b0), .COMP_OUT(na1435_3_i) );
// C_MULTFb//O_O2//      x40y52     80'h00_0018_13_A477_3EA6_0CCC
C_MULTFb   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1436_1 ( .COUTX(na1436_3), .COUTY1(na1436_4), .COUTY2(na1436_5), .POUTY1(na1436_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1415_3), .CINY1(na1435_4),
                      .CINY2(na1435_5), .PINX(1'b0), .PINY1(na1435_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_O2/AND/      x40y53     80'h00_0078_35_A471_3C88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1437_1 ( .OUT(na1437_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1436_4), .PINX(1'b0), .PINY1(na1436_7) );
C_O_O2     #(.CPE_CFG ()) 
           _a1437_3 ( .COMP_OUT(na1437_3_i), .COMB1(1'b0), .COMB2(na1437_2) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1437_4 ( .OUT(na1437_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1436_4), .PINX(1'b0), .PINY1(na1436_7) );
C_CPlines  #(.CPE_CFG (19'h3_5A47)) 
           _a1437_6 ( .COUTX(na1437_3), .COUTY1(na1437_4), .COUTY2(na1437_5), .POUTY1(na1437_7), .POUTY2(na1437_8), .CINX(1'b0), .CINY1(na1436_4),
                      .CINY2(na1436_5), .PINX(1'b0), .PINY1(na1436_7), .PINY2(1'b0), .OUT1(na1437_1), .OUT2(na1437_2), .COMP_OUT(na1437_3_i) );
// C_MULT///MULT/      x40y54     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1438_1 ( .COUTY1(na1438_4), .COUTY2(na1438_5), .POUTY1(na1438_7), .POUTY2(na1438_8), .IN1(~na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1417_3),
                      .CINY1(na1437_4), .CINY2(na1437_5), .PINX(na1417_6), .PINY1(na1437_7), .PINY2(na1437_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y55     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1439_1 ( .COUTX(na1439_3), .COUTY1(na1439_4), .COUTY2(na1439_5), .POUTX(na1439_6), .POUTY1(na1439_7), .POUTY2(na1439_8),
                      .IN1(na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1418_3), .CINY1(na1438_4), .CINY2(na1438_5), .PINX(na1418_6), .PINY1(na1438_7), .PINY2(na1438_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1440_1 ( .COUTX(na1440_3), .COUTY1(na1440_4), .COUTY2(na1440_5), .POUTX(na1440_6), .POUTY1(na1440_7), .POUTY2(na1440_8),
                      .IN1(~na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1419_3), .CINY1(na1439_4), .CINY2(na1439_5), .PINX(na1419_6), .PINY1(na1439_7), .PINY2(na1439_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1441_1 ( .COUTX(na1441_3), .COUTY1(na1441_4), .COUTY2(na1441_5), .POUTX(na1441_6), .POUTY1(na1441_7), .POUTY2(na1441_8),
                      .IN1(na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1420_3), .CINY1(na1440_4), .CINY2(na1440_5), .PINX(na1420_6), .PINY1(na1440_7), .PINY2(na1440_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1442_1 ( .COUTX(na1442_3), .COUTY1(na1442_4), .COUTY2(na1442_5), .POUTX(na1442_6), .POUTY1(na1442_7), .POUTY2(na1442_8),
                      .IN1(~na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1421_3), .CINY1(na1441_4), .CINY2(na1441_5), .PINX(na1421_6), .PINY1(na1441_7), .PINY2(na1441_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1443_1 ( .COUTX(na1443_3), .COUTY1(na1443_4), .COUTY2(na1443_5), .POUTX(na1443_6), .POUTY1(na1443_7), .POUTY2(na1443_8),
                      .IN1(na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1422_3), .CINY1(na1442_4), .CINY2(na1442_5), .PINX(na1422_6), .PINY1(na1442_7), .PINY2(na1442_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1444_1 ( .COUTX(na1444_3), .COUTY1(na1444_4), .COUTY2(na1444_5), .POUTX(na1444_6), .POUTY1(na1444_7), .POUTY2(na1444_8),
                      .IN1(~na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1423_3), .CINY1(na1443_4), .CINY2(na1443_5), .PINX(na1423_6), .PINY1(na1443_7), .PINY2(na1443_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y61     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1445_1 ( .COUTX(na1445_3), .COUTY1(na1445_4), .COUTY2(na1445_5), .POUTX(na1445_6), .POUTY1(na1445_7), .POUTY2(na1445_8),
                      .IN1(na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1424_3), .CINY1(na1444_4), .CINY2(na1444_5), .PINX(na1424_6), .PINY1(na1444_7), .PINY2(na1444_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y62     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1446_1 ( .COUTX(na1446_3), .COUTY1(na1446_4), .COUTY2(na1446_5), .POUTX(na1446_6), .POUTY1(na1446_7), .POUTY2(na1446_8),
                      .IN1(~na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1425_3), .CINY1(na1445_4), .CINY2(na1445_5), .PINX(na1425_6), .PINY1(na1445_7), .PINY2(na1445_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y63     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1447_1 ( .COUTX(na1447_3), .COUTY1(na1447_4), .COUTY2(na1447_5), .POUTX(na1447_6), .POUTY1(na1447_7), .POUTY2(na1447_8),
                      .IN1(na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1426_3), .CINY1(na1446_4), .CINY2(na1446_5), .PINX(na1426_6), .PINY1(na1446_7), .PINY2(na1446_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y64     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1448_1 ( .COUTX(na1448_3), .COUTY1(na1448_4), .COUTY2(na1448_5), .POUTX(na1448_6), .POUTY1(na1448_7), .POUTY2(na1448_8),
                      .IN1(~na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1427_3), .CINY1(na1447_4), .CINY2(na1447_5), .PINX(na1427_6), .PINY1(na1447_7), .PINY2(na1447_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y65     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1449_1 ( .COUTX(na1449_3), .COUTY1(na1449_4), .COUTY2(na1449_5), .POUTX(na1449_6), .POUTY1(na1449_7), .POUTY2(na1449_8),
                      .IN1(na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1428_3), .CINY1(na1448_4), .CINY2(na1448_5), .PINX(na1428_6), .PINY1(na1448_7), .PINY2(na1448_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y66     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1450_1 ( .COUTX(na1450_3), .COUTY1(na1450_4), .COUTY2(na1450_5), .POUTX(na1450_6), .POUTY1(na1450_7), .POUTY2(na1450_8),
                      .IN1(~na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1429_3), .CINY1(na1449_4), .CINY2(na1449_5), .PINX(na1429_6), .PINY1(na1449_7), .PINY2(na1449_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y67     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1451_1 ( .COUTX(na1451_3), .COUTY1(na1451_4), .COUTY2(na1451_5), .POUTX(na1451_6), .POUTY1(na1451_7), .POUTY2(na1451_8),
                      .IN1(na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1430_3), .CINY1(na1450_4), .CINY2(na1450_5), .PINX(na1430_6), .PINY1(na1450_7), .PINY2(na1450_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y68     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1452_1 ( .COUTX(na1452_3), .COUTY1(na1452_4), .COUTY2(na1452_5), .POUTX(na1452_6), .POUTY1(na1452_7), .POUTY2(na1452_8),
                      .IN1(~na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1431_3), .CINY1(na1451_4), .CINY2(na1451_5), .PINX(na1431_6), .PINY1(na1451_7), .PINY2(na1451_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y69     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1453_1 ( .COUTX(na1453_3), .COUTY1(na1453_4), .COUTY2(na1453_5), .POUTX(na1453_6), .POUTY1(na1453_7), .POUTY2(na1453_8),
                      .IN1(na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1432_3), .CINY1(na1452_4), .CINY2(na1452_5), .PINX(na1432_6), .PINY1(na1452_7), .PINY2(na1452_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x40y70     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1454_1 ( .COUTX(na1454_3), .COUTY1(na1454_4), .COUTY2(na1454_5), .POUTX(na1454_6), .POUTY1(na1454_7), .POUTY2(na1454_8),
                      .IN1(~na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1433_3), .CINY1(na1453_4), .CINY2(na1453_5), .PINX(na1433_6), .PINY1(na1453_7), .PINY2(na1453_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x40y71     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1455_3 ( .COMP_OUT(na1455_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1455_4 ( .OUT(na1455_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1454_4), .PINX(1'b0), .PINY1(na1454_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1455_6 ( .COUTX(na1455_3), .POUTX(na1455_6), .CINX(1'b0), .CINY1(na1454_4), .CINY2(na1454_5), .PINX(1'b0), .PINY1(na1454_7),
                      .PINY2(na1454_8), .OUT1(1'b0), .OUT2(na1455_2), .COMP_OUT(na1455_3_i) );
// C_AND///AND/      x41y51     80'h00_0078_12_0000_0C88_F0F0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1456_1 ( .OUT(na1456_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1456_4 ( .OUT(na1456_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1456_6 ( .COUTY1(na1456_4), .POUTY1(na1456_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1456_1), .OUT2(na1456_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x41y52     80'h00_0018_04_2056_5888_0CCF
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1457_1 ( .OUT(na1457_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(na1436_3), .CINY1(na1456_4), .PINX(1'b0), .PINY1(na1456_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1457_3 ( .COMP_OUT(na1457_3_i), .COMB1(na1457_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1457_6 ( .COUTY1(na1457_4), .COUTY2(na1457_5), .POUTY1(na1457_7), .CINX(na1436_3), .CINY1(na1456_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1456_7), .PINY2(1'b0), .OUT1(na1457_1), .OUT2(1'b0), .COMP_OUT(na1457_3_i) );
// C_MULTFa//O_O2//      x41y53     80'h00_0018_13_A477_34A6_0CCC
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1458_1 ( .COUTX(na1458_3), .COUTY1(na1458_4), .COUTY2(na1458_5), .POUTY1(na1458_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1437_3), .CINY1(na1457_4),
                      .CINY2(na1457_5), .PINX(1'b0), .PINY1(na1457_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x41y54     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1459_1 ( .OUT(na1459_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1458_4), .PINX(1'b0), .PINY1(na1458_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1459_3 ( .COMP_OUT(na1459_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1459_4 ( .OUT(na1459_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1458_4), .PINX(1'b0), .PINY1(na1458_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1459_6 ( .COUTX(na1459_3), .COUTY1(na1459_4), .COUTY2(na1459_5), .POUTY1(na1459_7), .POUTY2(na1459_8), .CINX(1'b0), .CINY1(na1458_4),
                      .CINY2(na1458_5), .PINX(1'b0), .PINY1(na1458_7), .PINY2(1'b0), .OUT1(na1459_1), .OUT2(na1459_2), .COMP_OUT(na1459_3_i) );
// C_MULT///MULT/      x41y55     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1460_1 ( .COUTY1(na1460_4), .COUTY2(na1460_5), .POUTY1(na1460_7), .POUTY2(na1460_8), .IN1(na1131_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1130_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1439_3),
                      .CINY1(na1459_4), .CINY2(na1459_5), .PINX(na1439_6), .PINY1(na1459_7), .PINY2(na1459_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y56     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1461_1 ( .COUTX(na1461_3), .COUTY1(na1461_4), .COUTY2(na1461_5), .POUTX(na1461_6), .POUTY1(na1461_7), .POUTY2(na1461_8),
                      .IN1(~na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1440_3), .CINY1(na1460_4), .CINY2(na1460_5), .PINX(na1440_6), .PINY1(na1460_7), .PINY2(na1460_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1462_1 ( .COUTX(na1462_3), .COUTY1(na1462_4), .COUTY2(na1462_5), .POUTX(na1462_6), .POUTY1(na1462_7), .POUTY2(na1462_8),
                      .IN1(na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1441_3), .CINY1(na1461_4), .CINY2(na1461_5), .PINX(na1441_6), .PINY1(na1461_7), .PINY2(na1461_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1463_1 ( .COUTX(na1463_3), .COUTY1(na1463_4), .COUTY2(na1463_5), .POUTX(na1463_6), .POUTY1(na1463_7), .POUTY2(na1463_8),
                      .IN1(~na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1442_3), .CINY1(na1462_4), .CINY2(na1462_5), .PINX(na1442_6), .PINY1(na1462_7), .PINY2(na1462_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1464_1 ( .COUTX(na1464_3), .COUTY1(na1464_4), .COUTY2(na1464_5), .POUTX(na1464_6), .POUTY1(na1464_7), .POUTY2(na1464_8),
                      .IN1(na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1443_3), .CINY1(na1463_4), .CINY2(na1463_5), .PINX(na1443_6), .PINY1(na1463_7), .PINY2(na1463_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1465_1 ( .COUTX(na1465_3), .COUTY1(na1465_4), .COUTY2(na1465_5), .POUTX(na1465_6), .POUTY1(na1465_7), .POUTY2(na1465_8),
                      .IN1(~na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1444_3), .CINY1(na1464_4), .CINY2(na1464_5), .PINX(na1444_6), .PINY1(na1464_7), .PINY2(na1464_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y61     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1466_1 ( .COUTX(na1466_3), .COUTY1(na1466_4), .COUTY2(na1466_5), .POUTX(na1466_6), .POUTY1(na1466_7), .POUTY2(na1466_8),
                      .IN1(na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1445_3), .CINY1(na1465_4), .CINY2(na1465_5), .PINX(na1445_6), .PINY1(na1465_7), .PINY2(na1465_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y62     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1467_1 ( .COUTX(na1467_3), .COUTY1(na1467_4), .COUTY2(na1467_5), .POUTX(na1467_6), .POUTY1(na1467_7), .POUTY2(na1467_8),
                      .IN1(~na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1446_3), .CINY1(na1466_4), .CINY2(na1466_5), .PINX(na1446_6), .PINY1(na1466_7), .PINY2(na1466_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y63     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1468_1 ( .COUTX(na1468_3), .COUTY1(na1468_4), .COUTY2(na1468_5), .POUTX(na1468_6), .POUTY1(na1468_7), .POUTY2(na1468_8),
                      .IN1(na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1447_3), .CINY1(na1467_4), .CINY2(na1467_5), .PINX(na1447_6), .PINY1(na1467_7), .PINY2(na1467_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y64     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1469_1 ( .COUTX(na1469_3), .COUTY1(na1469_4), .COUTY2(na1469_5), .POUTX(na1469_6), .POUTY1(na1469_7), .POUTY2(na1469_8),
                      .IN1(~na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1448_3), .CINY1(na1468_4), .CINY2(na1468_5), .PINX(na1448_6), .PINY1(na1468_7), .PINY2(na1468_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y65     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1470_1 ( .COUTX(na1470_3), .COUTY1(na1470_4), .COUTY2(na1470_5), .POUTX(na1470_6), .POUTY1(na1470_7), .POUTY2(na1470_8),
                      .IN1(na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1449_3), .CINY1(na1469_4), .CINY2(na1469_5), .PINX(na1449_6), .PINY1(na1469_7), .PINY2(na1469_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y66     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1471_1 ( .COUTX(na1471_3), .COUTY1(na1471_4), .COUTY2(na1471_5), .POUTX(na1471_6), .POUTY1(na1471_7), .POUTY2(na1471_8),
                      .IN1(~na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1450_3), .CINY1(na1470_4), .CINY2(na1470_5), .PINX(na1450_6), .PINY1(na1470_7), .PINY2(na1470_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y67     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1472_1 ( .COUTX(na1472_3), .COUTY1(na1472_4), .COUTY2(na1472_5), .POUTX(na1472_6), .POUTY1(na1472_7), .POUTY2(na1472_8),
                      .IN1(na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1451_3), .CINY1(na1471_4), .CINY2(na1471_5), .PINX(na1451_6), .PINY1(na1471_7), .PINY2(na1471_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y68     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1473_1 ( .COUTX(na1473_3), .COUTY1(na1473_4), .COUTY2(na1473_5), .POUTX(na1473_6), .POUTY1(na1473_7), .POUTY2(na1473_8),
                      .IN1(~na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1452_3), .CINY1(na1472_4), .CINY2(na1472_5), .PINX(na1452_6), .PINY1(na1472_7), .PINY2(na1472_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y69     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1474_1 ( .COUTX(na1474_3), .COUTY1(na1474_4), .COUTY2(na1474_5), .POUTX(na1474_6), .POUTY1(na1474_7), .POUTY2(na1474_8),
                      .IN1(na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1453_3), .CINY1(na1473_4), .CINY2(na1473_5), .PINX(na1453_6), .PINY1(na1473_7), .PINY2(na1473_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y70     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1475_1 ( .COUTX(na1475_3), .COUTY1(na1475_4), .COUTY2(na1475_5), .POUTX(na1475_6), .POUTY1(na1475_7), .POUTY2(na1475_8),
                      .IN1(~na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1454_3), .CINY1(na1474_4), .CINY2(na1474_5), .PINX(na1454_6), .PINY1(na1474_7), .PINY2(na1474_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x41y71     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1476_1 ( .COUTX(na1476_3), .COUTY1(na1476_4), .COUTY2(na1476_5), .POUTX(na1476_6), .POUTY1(na1476_7), .POUTY2(na1476_8),
                      .IN1(na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1455_3), .CINY1(na1475_4), .CINY2(na1475_5), .PINX(na1455_6), .PINY1(na1475_7), .PINY2(na1475_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x41y72     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1477_3 ( .COMP_OUT(na1477_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1477_4 ( .OUT(na1477_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1476_4), .PINX(1'b0), .PINY1(na1476_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1477_6 ( .COUTX(na1477_3), .POUTX(na1477_6), .CINX(1'b0), .CINY1(na1476_4), .CINY2(na1476_5), .PINX(1'b0), .PINY1(na1476_7),
                      .PINY2(na1476_8), .OUT1(1'b0), .OUT2(na1477_2), .COMP_OUT(na1477_3_i) );
// C_AND///AND/      x42y52     80'h00_0078_12_0000_0C88_FFF0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1478_1 ( .OUT(na1478_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1478_4 ( .OUT(na1478_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1478_6 ( .COUTY1(na1478_4), .POUTY1(na1478_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1478_1), .OUT2(na1478_2), .COMP_OUT(1'b0) );
// C_OR//O_O1//      x42y53     80'h00_0018_04_2056_5EEE_0CC0
C_OR       #(.CPE_CFG (9'b0_0001_0110)) 
           _a1479_1 ( .OUT(na1479_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(na1458_3), .CINY1(na1478_4), .PINX(1'b0), .PINY1(na1478_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1479_3 ( .COMP_OUT(na1479_3_i), .COMB1(na1479_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1479_6 ( .COUTY1(na1479_4), .COUTY2(na1479_5), .POUTY1(na1479_7), .CINX(na1458_3), .CINY1(na1478_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1478_7), .PINY2(1'b0), .OUT1(na1479_1), .OUT2(1'b0), .COMP_OUT(na1479_3_i) );
// C_MULTFb//O_O2//      x42y54     80'h00_0018_13_A477_3EA6_0CCC
C_MULTFb   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1480_1 ( .COUTX(na1480_3), .COUTY1(na1480_4), .COUTY2(na1480_5), .POUTY1(na1480_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1459_3), .CINY1(na1479_4),
                      .CINY2(na1479_5), .PINX(1'b0), .PINY1(na1479_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_O2/AND/      x42y55     80'h00_0078_35_A471_3C88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1481_1 ( .OUT(na1481_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1480_4), .PINX(1'b0), .PINY1(na1480_7) );
C_O_O2     #(.CPE_CFG ()) 
           _a1481_3 ( .COMP_OUT(na1481_3_i), .COMB1(1'b0), .COMB2(na1481_2) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1481_4 ( .OUT(na1481_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1480_4), .PINX(1'b0), .PINY1(na1480_7) );
C_CPlines  #(.CPE_CFG (19'h3_5A47)) 
           _a1481_6 ( .COUTX(na1481_3), .COUTY1(na1481_4), .COUTY2(na1481_5), .POUTY1(na1481_7), .POUTY2(na1481_8), .CINX(1'b0), .CINY1(na1480_4),
                      .CINY2(na1480_5), .PINX(1'b0), .PINY1(na1480_7), .PINY2(1'b0), .OUT1(na1481_1), .OUT2(na1481_2), .COMP_OUT(na1481_3_i) );
// C_MULT///MULT/      x42y56     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1482_1 ( .OUT1(na1482_1), .OUT2(na1482_2), .COUTY1(na1482_4), .COUTY2(na1482_5), .POUTY1(na1482_7), .POUTY2(na1482_8), .IN1(~na1131_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1130_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1461_3), .CINY1(na1481_4), .CINY2(na1481_5), .PINX(na1461_6), .PINY1(na1481_7), .PINY2(na1481_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y57     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1483_1 ( .COUTX(na1483_3), .COUTY1(na1483_4), .COUTY2(na1483_5), .POUTX(na1483_6), .POUTY1(na1483_7), .POUTY2(na1483_8),
                      .IN1(na1132_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1131_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1462_3), .CINY1(na1482_4), .CINY2(na1482_5), .PINX(na1462_6), .PINY1(na1482_7), .PINY2(na1482_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y58     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1484_1 ( .COUTX(na1484_3), .COUTY1(na1484_4), .COUTY2(na1484_5), .POUTX(na1484_6), .POUTY1(na1484_7), .POUTY2(na1484_8),
                      .IN1(~na1133_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1132_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1463_3), .CINY1(na1483_4), .CINY2(na1483_5), .PINX(na1463_6), .PINY1(na1483_7), .PINY2(na1483_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y59     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1485_1 ( .COUTX(na1485_3), .COUTY1(na1485_4), .COUTY2(na1485_5), .POUTX(na1485_6), .POUTY1(na1485_7), .POUTY2(na1485_8),
                      .IN1(na1134_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1133_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1464_3), .CINY1(na1484_4), .CINY2(na1484_5), .PINX(na1464_6), .PINY1(na1484_7), .PINY2(na1484_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y60     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1486_1 ( .COUTX(na1486_3), .COUTY1(na1486_4), .COUTY2(na1486_5), .POUTX(na1486_6), .POUTY1(na1486_7), .POUTY2(na1486_8),
                      .IN1(~na1135_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1134_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1465_3), .CINY1(na1485_4), .CINY2(na1485_5), .PINX(na1465_6), .PINY1(na1485_7), .PINY2(na1485_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y61     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1487_1 ( .COUTX(na1487_3), .COUTY1(na1487_4), .COUTY2(na1487_5), .POUTX(na1487_6), .POUTY1(na1487_7), .POUTY2(na1487_8),
                      .IN1(na1136_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1135_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1466_3), .CINY1(na1486_4), .CINY2(na1486_5), .PINX(na1466_6), .PINY1(na1486_7), .PINY2(na1486_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y62     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1488_1 ( .COUTX(na1488_3), .COUTY1(na1488_4), .COUTY2(na1488_5), .POUTX(na1488_6), .POUTY1(na1488_7), .POUTY2(na1488_8),
                      .IN1(~na1137_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1136_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1467_3), .CINY1(na1487_4), .CINY2(na1487_5), .PINX(na1467_6), .PINY1(na1487_7), .PINY2(na1487_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y63     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1489_1 ( .COUTX(na1489_3), .COUTY1(na1489_4), .COUTY2(na1489_5), .POUTX(na1489_6), .POUTY1(na1489_7), .POUTY2(na1489_8),
                      .IN1(na1138_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1137_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1468_3), .CINY1(na1488_4), .CINY2(na1488_5), .PINX(na1468_6), .PINY1(na1488_7), .PINY2(na1488_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y64     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1490_1 ( .COUTX(na1490_3), .COUTY1(na1490_4), .COUTY2(na1490_5), .POUTX(na1490_6), .POUTY1(na1490_7), .POUTY2(na1490_8),
                      .IN1(~na1139_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1138_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1469_3), .CINY1(na1489_4), .CINY2(na1489_5), .PINX(na1469_6), .PINY1(na1489_7), .PINY2(na1489_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y65     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1491_1 ( .COUTX(na1491_3), .COUTY1(na1491_4), .COUTY2(na1491_5), .POUTX(na1491_6), .POUTY1(na1491_7), .POUTY2(na1491_8),
                      .IN1(na1140_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1139_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1470_3), .CINY1(na1490_4), .CINY2(na1490_5), .PINX(na1470_6), .PINY1(na1490_7), .PINY2(na1490_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y66     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1492_1 ( .COUTX(na1492_3), .COUTY1(na1492_4), .COUTY2(na1492_5), .POUTX(na1492_6), .POUTY1(na1492_7), .POUTY2(na1492_8),
                      .IN1(~na1141_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1140_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1471_3), .CINY1(na1491_4), .CINY2(na1491_5), .PINX(na1471_6), .PINY1(na1491_7), .PINY2(na1491_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y67     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1493_1 ( .COUTX(na1493_3), .COUTY1(na1493_4), .COUTY2(na1493_5), .POUTX(na1493_6), .POUTY1(na1493_7), .POUTY2(na1493_8),
                      .IN1(na1142_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1141_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1472_3), .CINY1(na1492_4), .CINY2(na1492_5), .PINX(na1472_6), .PINY1(na1492_7), .PINY2(na1492_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y68     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1494_1 ( .COUTX(na1494_3), .COUTY1(na1494_4), .COUTY2(na1494_5), .POUTX(na1494_6), .POUTY1(na1494_7), .POUTY2(na1494_8),
                      .IN1(~na1143_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1142_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1473_3), .CINY1(na1493_4), .CINY2(na1493_5), .PINX(na1473_6), .PINY1(na1493_7), .PINY2(na1493_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y69     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1495_1 ( .COUTX(na1495_3), .COUTY1(na1495_4), .COUTY2(na1495_5), .POUTX(na1495_6), .POUTY1(na1495_7), .POUTY2(na1495_8),
                      .IN1(na1144_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1143_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1474_3), .CINY1(na1494_4), .CINY2(na1494_5), .PINX(na1474_6), .PINY1(na1494_7), .PINY2(na1494_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y70     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1496_1 ( .COUTX(na1496_3), .COUTY1(na1496_4), .COUTY2(na1496_5), .POUTX(na1496_6), .POUTY1(na1496_7), .POUTY2(na1496_8),
                      .IN1(~na1145_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1144_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1475_3), .CINY1(na1495_4), .CINY2(na1495_5), .PINX(na1475_6), .PINY1(na1495_7), .PINY2(na1495_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y71     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1497_1 ( .COUTX(na1497_3), .COUTY1(na1497_4), .COUTY2(na1497_5), .POUTX(na1497_6), .POUTY1(na1497_7), .POUTY2(na1497_8),
                      .IN1(na1146_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1145_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1476_3), .CINY1(na1496_4), .CINY2(na1496_5), .PINX(na1476_6), .PINY1(na1496_7), .PINY2(na1496_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x42y72     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1498_1 ( .COUTX(na1498_3), .COUTY1(na1498_4), .COUTY2(na1498_5), .POUTX(na1498_6), .POUTY1(na1498_7), .POUTY2(na1498_8),
                      .IN1(~na1147_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1146_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1477_3), .CINY1(na1497_4), .CINY2(na1497_5), .PINX(na1477_6), .PINY1(na1497_7), .PINY2(na1497_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x42y73     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1499_3 ( .COMP_OUT(na1499_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1499_4 ( .OUT(na1499_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1498_4), .PINX(1'b0), .PINY1(na1498_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1499_6 ( .COUTX(na1499_3), .POUTX(na1499_6), .CINX(1'b0), .CINY1(na1498_4), .CINY2(na1498_5), .PINX(1'b0), .PINY1(na1498_7),
                      .PINY2(na1498_8), .OUT1(1'b0), .OUT2(na1499_2), .COMP_OUT(na1499_3_i) );
// C_AND///AND/      x43y53     80'h00_0078_12_0000_0C88_F0F0
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1500_1 ( .OUT(na1500_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1500_4 ( .OUT(na1500_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1500_6 ( .COUTY1(na1500_4), .POUTY1(na1500_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1500_1), .OUT2(na1500_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x43y54     80'h00_0018_04_2056_5888_0CCF
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1501_1 ( .OUT(na1501_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(na1480_3), .CINY1(na1500_4), .PINX(1'b0), .PINY1(na1500_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1501_3 ( .COMP_OUT(na1501_3_i), .COMB1(na1501_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1501_6 ( .COUTY1(na1501_4), .COUTY2(na1501_5), .POUTY1(na1501_7), .CINX(na1480_3), .CINY1(na1500_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1500_7), .PINY2(1'b0), .OUT1(na1501_1), .OUT2(1'b0), .COMP_OUT(na1501_3_i) );
// C_MULTFa//O_O2//      x43y55     80'h00_0018_13_A477_34A6_0CCC
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1502_1 ( .COUTY1(na1502_4), .COUTY2(na1502_5), .POUTY1(na1502_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1),
                      .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1481_3), .CINY1(na1501_4), .CINY2(na1501_5),
                      .PINX(1'b0), .PINY1(na1501_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x43y56     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1503_1 ( .OUT(na1503_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1502_4), .PINX(1'b0), .PINY1(na1502_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1503_3 ( .COMP_OUT(na1503_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1503_4 ( .OUT(na1503_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1502_4), .PINX(1'b0), .PINY1(na1502_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1503_6 ( .COUTY1(na1503_4), .COUTY2(na1503_5), .POUTY1(na1503_7), .POUTY2(na1503_8), .CINX(1'b0), .CINY1(na1502_4), .CINY2(na1502_5),
                      .PINX(1'b0), .PINY1(na1502_7), .PINY2(1'b0), .OUT1(na1503_1), .OUT2(na1503_2), .COMP_OUT(na1503_3_i) );
// C_MULT///MULT/      x43y57     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1504_1 ( .OUT1(na1504_1), .OUT2(na1504_2), .COUTY1(na1504_4), .COUTY2(na1504_5), .POUTY1(na1504_7), .POUTY2(na1504_8), .IN1(na1131_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1131_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1130_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1483_3), .CINY1(na1503_4), .CINY2(na1503_5), .PINX(na1483_6), .PINY1(na1503_7), .PINY2(na1503_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y58     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1505_1 ( .OUT1(na1505_1), .OUT2(na1505_2), .COUTY1(na1505_4), .COUTY2(na1505_5), .POUTY1(na1505_7), .POUTY2(na1505_8), .IN1(~na1132_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1132_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1131_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1484_3), .CINY1(na1504_4), .CINY2(na1504_5), .PINX(na1484_6), .PINY1(na1504_7), .PINY2(na1504_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y59     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1506_1 ( .OUT1(na1506_1), .OUT2(na1506_2), .COUTY1(na1506_4), .COUTY2(na1506_5), .POUTY1(na1506_7), .POUTY2(na1506_8), .IN1(na1133_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1133_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1132_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1485_3), .CINY1(na1505_4), .CINY2(na1505_5), .PINX(na1485_6), .PINY1(na1505_7), .PINY2(na1505_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y60     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1507_1 ( .OUT1(na1507_1), .OUT2(na1507_2), .COUTY1(na1507_4), .COUTY2(na1507_5), .POUTY1(na1507_7), .POUTY2(na1507_8), .IN1(~na1134_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1134_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1133_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1486_3), .CINY1(na1506_4), .CINY2(na1506_5), .PINX(na1486_6), .PINY1(na1506_7), .PINY2(na1506_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y61     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1508_1 ( .OUT1(na1508_1), .OUT2(na1508_2), .COUTY1(na1508_4), .COUTY2(na1508_5), .POUTY1(na1508_7), .POUTY2(na1508_8), .IN1(na1135_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1135_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1134_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1487_3), .CINY1(na1507_4), .CINY2(na1507_5), .PINX(na1487_6), .PINY1(na1507_7), .PINY2(na1507_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y62     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1509_1 ( .OUT1(na1509_1), .OUT2(na1509_2), .COUTY1(na1509_4), .COUTY2(na1509_5), .POUTY1(na1509_7), .POUTY2(na1509_8), .IN1(~na1136_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1136_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1135_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1488_3), .CINY1(na1508_4), .CINY2(na1508_5), .PINX(na1488_6), .PINY1(na1508_7), .PINY2(na1508_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y63     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1510_1 ( .OUT1(na1510_1), .OUT2(na1510_2), .COUTY1(na1510_4), .COUTY2(na1510_5), .POUTY1(na1510_7), .POUTY2(na1510_8), .IN1(na1137_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1137_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1136_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1489_3), .CINY1(na1509_4), .CINY2(na1509_5), .PINX(na1489_6), .PINY1(na1509_7), .PINY2(na1509_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y64     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1511_1 ( .OUT1(na1511_1), .OUT2(na1511_2), .COUTY1(na1511_4), .COUTY2(na1511_5), .POUTY1(na1511_7), .POUTY2(na1511_8), .IN1(~na1138_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1138_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1137_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1490_3), .CINY1(na1510_4), .CINY2(na1510_5), .PINX(na1490_6), .PINY1(na1510_7), .PINY2(na1510_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y65     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1512_1 ( .OUT1(na1512_1), .OUT2(na1512_2), .COUTY1(na1512_4), .COUTY2(na1512_5), .POUTY1(na1512_7), .POUTY2(na1512_8), .IN1(na1139_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1139_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1138_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1491_3), .CINY1(na1511_4), .CINY2(na1511_5), .PINX(na1491_6), .PINY1(na1511_7), .PINY2(na1511_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y66     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1513_1 ( .OUT1(na1513_1), .OUT2(na1513_2), .COUTY1(na1513_4), .COUTY2(na1513_5), .POUTY1(na1513_7), .POUTY2(na1513_8), .IN1(~na1140_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1140_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1139_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1492_3), .CINY1(na1512_4), .CINY2(na1512_5), .PINX(na1492_6), .PINY1(na1512_7), .PINY2(na1512_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y67     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1514_1 ( .OUT1(na1514_1), .OUT2(na1514_2), .COUTY1(na1514_4), .COUTY2(na1514_5), .POUTY1(na1514_7), .POUTY2(na1514_8), .IN1(na1141_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1141_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1140_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1493_3), .CINY1(na1513_4), .CINY2(na1513_5), .PINX(na1493_6), .PINY1(na1513_7), .PINY2(na1513_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y68     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1515_1 ( .OUT1(na1515_1), .OUT2(na1515_2), .COUTY1(na1515_4), .COUTY2(na1515_5), .POUTY1(na1515_7), .POUTY2(na1515_8), .IN1(~na1142_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1142_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1141_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1494_3), .CINY1(na1514_4), .CINY2(na1514_5), .PINX(na1494_6), .PINY1(na1514_7), .PINY2(na1514_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y69     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1516_1 ( .OUT1(na1516_1), .OUT2(na1516_2), .COUTY1(na1516_4), .COUTY2(na1516_5), .POUTY1(na1516_7), .POUTY2(na1516_8), .IN1(na1143_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1143_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1142_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1495_3), .CINY1(na1515_4), .CINY2(na1515_5), .PINX(na1495_6), .PINY1(na1515_7), .PINY2(na1515_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y70     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1517_1 ( .COUTY1(na1517_4), .COUTY2(na1517_5), .POUTY1(na1517_7), .POUTY2(na1517_8), .IN1(~na1144_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na1144_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1143_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1496_3),
                      .CINY1(na1516_4), .CINY2(na1516_5), .PINX(na1496_6), .PINY1(na1516_7), .PINY2(na1516_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y71     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1518_1 ( .COUTY1(na1518_4), .COUTY2(na1518_5), .POUTY1(na1518_7), .POUTY2(na1518_8), .IN1(na1145_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1145_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1144_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1497_3),
                      .CINY1(na1517_4), .CINY2(na1517_5), .PINX(na1497_6), .PINY1(na1517_7), .PINY2(na1517_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y72     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1519_1 ( .COUTY1(na1519_4), .COUTY2(na1519_5), .POUTY1(na1519_7), .POUTY2(na1519_8), .IN1(~na1146_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na1146_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1145_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1498_3),
                      .CINY1(na1518_4), .CINY2(na1518_5), .PINX(na1498_6), .PINY1(na1518_7), .PINY2(na1518_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x43y73     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1520_1 ( .COUTY1(na1520_4), .COUTY2(na1520_5), .POUTY1(na1520_7), .POUTY2(na1520_8), .IN1(na1147_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1147_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1146_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1499_3),
                      .CINY1(na1519_4), .CINY2(na1519_5), .PINX(na1499_6), .PINY1(na1519_7), .PINY2(na1519_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x43y74     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1521_3 ( .COMP_OUT(na1521_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1521_4 ( .OUT(na1521_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1520_4), .PINX(1'b0), .PINY1(na1520_7) );
// C_///AND/      x45y73     80'h00_0060_00_0000_0C08_FFF0
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1522_4 ( .OUT(na1522_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
// C_AND//O_0/AND/      x45y74     80'h00_0078_09_6000_FC88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1523_1 ( .OUT(na1523_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na559_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a1523_3 ( .COMP_OUT(na1523_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1523_4 ( .OUT(na1523_2), .IN1(1'b1), .IN2(na559_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1523_6 ( .COUTX(na1523_3), .POUTX(na1523_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1523_1), .OUT2(na1523_2), .COMP_OUT(na1523_3_i) );
// C_AND//O_0/AND/      x45y75     80'h00_0078_09_6000_FC88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1524_1 ( .OUT(na1524_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na567_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a1524_3 ( .COMP_OUT(na1524_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1524_4 ( .OUT(na1524_2), .IN1(na567_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1524_6 ( .COUTX(na1524_3), .POUTX(na1524_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1524_1), .OUT2(na1524_2), .COMP_OUT(na1524_3_i) );
// C_AND//O_0/AND/      x45y76     80'h00_0078_09_6000_FC88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1525_1 ( .OUT(na1525_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na569_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a1525_3 ( .COMP_OUT(na1525_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1525_4 ( .OUT(na1525_2), .IN1(1'b1), .IN2(na569_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1525_6 ( .COUTX(na1525_3), .POUTX(na1525_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1525_1), .OUT2(na1525_2), .COMP_OUT(na1525_3_i) );
// C_AND//O_0/AND/      x45y77     80'h00_0078_09_6000_FC88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1526_1 ( .OUT(na1526_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na571_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a1526_3 ( .COMP_OUT(na1526_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1526_4 ( .OUT(na1526_2), .IN1(na571_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1526_6 ( .COUTX(na1526_3), .POUTX(na1526_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1526_1), .OUT2(na1526_2), .COMP_OUT(na1526_3_i) );
// C_AND//O_0/AND/      x45y78     80'h00_0078_09_6000_FC88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1527_1 ( .OUT(na1527_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na573_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a1527_3 ( .COMP_OUT(na1527_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1527_4 ( .OUT(na1527_2), .IN1(1'b1), .IN2(na573_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1527_6 ( .COUTX(na1527_3), .POUTX(na1527_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1527_1), .OUT2(na1527_2), .COMP_OUT(na1527_3_i) );
// C_AND//O_0/AND/      x45y79     80'h00_0078_09_6000_FC88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1528_1 ( .OUT(na1528_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na560_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a1528_3 ( .COMP_OUT(na1528_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1528_4 ( .OUT(na1528_2), .IN1(na560_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1528_6 ( .COUTX(na1528_3), .POUTX(na1528_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1528_1), .OUT2(na1528_2), .COMP_OUT(na1528_3_i) );
// C_AND//O_0/AND/      x45y80     80'h00_0078_09_6000_FC88_FCFC
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1529_1 ( .OUT(na1529_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(na562_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a1529_3 ( .COMP_OUT(na1529_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1529_4 ( .OUT(na1529_2), .IN1(1'b1), .IN2(na562_2), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1529_6 ( .COUTX(na1529_3), .POUTX(na1529_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1529_1), .OUT2(na1529_2), .COMP_OUT(na1529_3_i) );
// C_AND//O_0/AND/      x45y81     80'h00_0078_09_6000_FC88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1530_1 ( .OUT(na1530_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na564_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a1530_3 ( .COMP_OUT(na1530_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1530_4 ( .OUT(na1530_2), .IN1(na564_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1530_6 ( .COUTX(na1530_3), .POUTX(na1530_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1530_1), .OUT2(na1530_2), .COMP_OUT(na1530_3_i) );
// C_AND//O_0/AND/      x45y82     80'h00_0078_09_6000_FC88_FAFA
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1531_1 ( .OUT(na1531_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na564_2), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_O_0      #(.CPE_CFG ()) 
           _a1531_3 ( .COMP_OUT(na1531_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1531_4 ( .OUT(na1531_2), .IN1(na564_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_9600)) 
           _a1531_6 ( .COUTX(na1531_3), .POUTX(na1531_6), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1531_1), .OUT2(na1531_2), .COMP_OUT(na1531_3_i) );
// C_AND///AND/      x46y70     80'h00_0078_12_0000_0C88_3FAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1532_1 ( .OUT(na1532_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(~na60_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1532_4 ( .OUT(na1532_2), .IN1(1'b1), .IN2(1'b1), .IN3(na61_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1532_6 ( .COUTY1(na1532_4), .POUTY1(na1532_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1532_1), .OUT2(na1532_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x46y71     80'h00_0018_04_2056_5888_0CC0
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1533_1 ( .OUT(na1533_1), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1532_4), .PINX(1'b0), .PINY1(na1532_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1533_3 ( .COMP_OUT(na1533_3_i), .COMB1(na1533_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1533_6 ( .COUTY1(na1533_4), .COUTY2(na1533_5), .POUTY1(na1533_7), .CINX(1'b0), .CINY1(na1532_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1532_7), .PINY2(1'b0), .OUT1(na1533_1), .OUT2(1'b0), .COMP_OUT(na1533_3_i) );
// C_MULTFa//O_O2//      x46y72     80'h00_0018_13_A477_34A6_0C0C
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1534_1 ( .COUTX(na1534_3), .COUTY1(na1534_4), .COUTY2(na1534_5), .POUTY1(na1534_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b0), .IN4(1'b0),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1533_4),
                      .CINY2(na1533_5), .PINX(1'b0), .PINY1(na1533_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x46y73     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1535_1 ( .OUT(na1535_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1534_4), .PINX(1'b0), .PINY1(na1534_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1535_3 ( .COMP_OUT(na1535_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1535_4 ( .OUT(na1535_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1534_4), .PINX(1'b0), .PINY1(na1534_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1535_6 ( .COUTX(na1535_3), .COUTY1(na1535_4), .COUTY2(na1535_5), .POUTY1(na1535_7), .POUTY2(na1535_8), .CINX(1'b0), .CINY1(na1534_4),
                      .CINY2(na1534_5), .PINX(1'b0), .PINY1(na1534_7), .PINY2(1'b0), .OUT1(na1535_1), .OUT2(na1535_2), .COMP_OUT(na1535_3_i) );
// C_MULT///MULT/      x46y74     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1536_1 ( .COUTY1(na1536_4), .COUTY2(na1536_5), .POUTY1(na1536_7), .POUTY2(na1536_8), .IN1(na1523_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1523_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1522_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(1'b0),
                      .CINY1(na1535_4), .CINY2(na1535_5), .PINX(1'b0), .PINY1(na1535_7), .PINY2(na1535_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x46y75     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1537_1 ( .COUTX(na1537_3), .COUTY1(na1537_4), .COUTY2(na1537_5), .POUTX(na1537_6), .POUTY1(na1537_7), .POUTY2(na1537_8),
                      .IN1(na1524_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1524_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1523_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1536_4), .CINY2(na1536_5), .PINX(1'b0), .PINY1(na1536_7), .PINY2(na1536_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x46y76     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1538_1 ( .COUTX(na1538_3), .COUTY1(na1538_4), .COUTY2(na1538_5), .POUTX(na1538_6), .POUTY1(na1538_7), .POUTY2(na1538_8),
                      .IN1(na1525_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1525_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1524_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1537_4), .CINY2(na1537_5), .PINX(1'b0), .PINY1(na1537_7), .PINY2(na1537_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x46y77     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1539_1 ( .COUTX(na1539_3), .COUTY1(na1539_4), .COUTY2(na1539_5), .POUTX(na1539_6), .POUTY1(na1539_7), .POUTY2(na1539_8),
                      .IN1(na1526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1526_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1525_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1538_4), .CINY2(na1538_5), .PINX(1'b0), .PINY1(na1538_7), .PINY2(na1538_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x46y78     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1540_1 ( .COUTX(na1540_3), .COUTY1(na1540_4), .COUTY2(na1540_5), .POUTX(na1540_6), .POUTY1(na1540_7), .POUTY2(na1540_8),
                      .IN1(na1527_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1527_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1526_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1539_4), .CINY2(na1539_5), .PINX(1'b0), .PINY1(na1539_7), .PINY2(na1539_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x46y79     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1541_1 ( .COUTX(na1541_3), .COUTY1(na1541_4), .COUTY2(na1541_5), .POUTX(na1541_6), .POUTY1(na1541_7), .POUTY2(na1541_8),
                      .IN1(na1528_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1528_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1527_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1540_4), .CINY2(na1540_5), .PINX(1'b0), .PINY1(na1540_7), .PINY2(na1540_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x46y80     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1542_1 ( .COUTX(na1542_3), .COUTY1(na1542_4), .COUTY2(na1542_5), .POUTX(na1542_6), .POUTY1(na1542_7), .POUTY2(na1542_8),
                      .IN1(na1529_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1529_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1528_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1541_4), .CINY2(na1541_5), .PINX(1'b0), .PINY1(na1541_7), .PINY2(na1541_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x46y81     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1543_1 ( .COUTX(na1543_3), .COUTY1(na1543_4), .COUTY2(na1543_5), .POUTX(na1543_6), .POUTY1(na1543_7), .POUTY2(na1543_8),
                      .IN1(na1530_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1530_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1529_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1542_4), .CINY2(na1542_5), .PINX(1'b0), .PINY1(na1542_7), .PINY2(na1542_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x46y82     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1544_1 ( .COUTX(na1544_3), .COUTY1(na1544_4), .COUTY2(na1544_5), .POUTX(na1544_6), .POUTY1(na1544_7), .POUTY2(na1544_8),
                      .IN1(na1531_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1531_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1530_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(1'b0), .CINY1(na1543_4), .CINY2(na1543_5), .PINX(1'b0), .PINY1(na1543_7), .PINY2(na1543_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x46y83     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1545_3 ( .COMP_OUT(na1545_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1545_4 ( .OUT(na1545_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1544_4), .PINX(1'b0), .PINY1(na1544_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1545_6 ( .COUTX(na1545_3), .POUTX(na1545_6), .CINX(1'b0), .CINY1(na1544_4), .CINY2(na1544_5), .PINX(1'b0), .PINY1(na1544_7),
                      .PINY2(na1544_8), .OUT1(1'b0), .OUT2(na1545_2), .COMP_OUT(na1545_3_i) );
// C_AND///AND/      x47y71     80'h00_0078_12_0000_0C88_CFAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1546_1 ( .OUT(na1546_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(na63_1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1546_4 ( .OUT(na1546_2), .IN1(1'b1), .IN2(1'b1), .IN3(na65_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1546_6 ( .COUTY1(na1546_4), .POUTY1(na1546_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1546_1), .OUT2(na1546_2), .COMP_OUT(1'b0) );
// C_OR//O_O1//      x47y72     80'h00_0018_04_2056_5EEE_0CC0
C_OR       #(.CPE_CFG (9'b0_0001_0110)) 
           _a1547_1 ( .OUT(na1547_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(na1534_3), .CINY1(na1546_4), .PINX(1'b0), .PINY1(na1546_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1547_3 ( .COMP_OUT(na1547_3_i), .COMB1(na1547_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1547_6 ( .COUTY1(na1547_4), .COUTY2(na1547_5), .POUTY1(na1547_7), .CINX(na1534_3), .CINY1(na1546_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1546_7), .PINY2(1'b0), .OUT1(na1547_1), .OUT2(1'b0), .COMP_OUT(na1547_3_i) );
// C_MULTFb//O_O2//      x47y73     80'h00_0018_13_A477_3EA6_0CCC
C_MULTFb   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1548_1 ( .COUTX(na1548_3), .COUTY1(na1548_4), .COUTY2(na1548_5), .POUTY1(na1548_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1535_3), .CINY1(na1547_4),
                      .CINY2(na1547_5), .PINX(1'b0), .PINY1(na1547_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_O2/AND/      x47y74     80'h00_0078_35_A471_3C88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1549_1 ( .OUT(na1549_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1548_4), .PINX(1'b0), .PINY1(na1548_7) );
C_O_O2     #(.CPE_CFG ()) 
           _a1549_3 ( .COMP_OUT(na1549_3_i), .COMB1(1'b0), .COMB2(na1549_2) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1549_4 ( .OUT(na1549_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1548_4), .PINX(1'b0), .PINY1(na1548_7) );
C_CPlines  #(.CPE_CFG (19'h3_5A47)) 
           _a1549_6 ( .COUTX(na1549_3), .COUTY1(na1549_4), .COUTY2(na1549_5), .POUTY1(na1549_7), .POUTY2(na1549_8), .CINX(1'b0), .CINY1(na1548_4),
                      .CINY2(na1548_5), .PINX(1'b0), .PINY1(na1548_7), .PINY2(1'b0), .OUT1(na1549_1), .OUT2(na1549_2), .COMP_OUT(na1549_3_i) );
// C_MULT///MULT/      x47y75     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1550_1 ( .COUTY1(na1550_4), .COUTY2(na1550_5), .POUTY1(na1550_7), .POUTY2(na1550_8), .IN1(~na1523_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(~na1523_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1522_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1537_3),
                      .CINY1(na1549_4), .CINY2(na1549_5), .PINX(na1537_6), .PINY1(na1549_7), .PINY2(na1549_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x47y76     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1551_1 ( .COUTX(na1551_3), .COUTY1(na1551_4), .COUTY2(na1551_5), .POUTX(na1551_6), .POUTY1(na1551_7), .POUTY2(na1551_8),
                      .IN1(~na1524_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1524_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1523_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1538_3), .CINY1(na1550_4), .CINY2(na1550_5), .PINX(na1538_6), .PINY1(na1550_7), .PINY2(na1550_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x47y77     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1552_1 ( .COUTX(na1552_3), .COUTY1(na1552_4), .COUTY2(na1552_5), .POUTX(na1552_6), .POUTY1(na1552_7), .POUTY2(na1552_8),
                      .IN1(~na1525_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1525_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1524_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1539_3), .CINY1(na1551_4), .CINY2(na1551_5), .PINX(na1539_6), .PINY1(na1551_7), .PINY2(na1551_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x47y78     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1553_1 ( .COUTX(na1553_3), .COUTY1(na1553_4), .COUTY2(na1553_5), .POUTX(na1553_6), .POUTY1(na1553_7), .POUTY2(na1553_8),
                      .IN1(~na1526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1526_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1525_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1540_3), .CINY1(na1552_4), .CINY2(na1552_5), .PINX(na1540_6), .PINY1(na1552_7), .PINY2(na1552_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x47y79     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1554_1 ( .COUTX(na1554_3), .COUTY1(na1554_4), .COUTY2(na1554_5), .POUTX(na1554_6), .POUTY1(na1554_7), .POUTY2(na1554_8),
                      .IN1(~na1527_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1527_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1526_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1541_3), .CINY1(na1553_4), .CINY2(na1553_5), .PINX(na1541_6), .PINY1(na1553_7), .PINY2(na1553_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x47y80     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1555_1 ( .COUTX(na1555_3), .COUTY1(na1555_4), .COUTY2(na1555_5), .POUTX(na1555_6), .POUTY1(na1555_7), .POUTY2(na1555_8),
                      .IN1(~na1528_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1528_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1527_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1542_3), .CINY1(na1554_4), .CINY2(na1554_5), .PINX(na1542_6), .PINY1(na1554_7), .PINY2(na1554_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x47y81     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1556_1 ( .COUTX(na1556_3), .COUTY1(na1556_4), .COUTY2(na1556_5), .POUTX(na1556_6), .POUTY1(na1556_7), .POUTY2(na1556_8),
                      .IN1(~na1529_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1529_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1528_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1543_3), .CINY1(na1555_4), .CINY2(na1555_5), .PINX(na1543_6), .PINY1(na1555_7), .PINY2(na1555_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x47y82     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1557_1 ( .COUTX(na1557_3), .COUTY1(na1557_4), .COUTY2(na1557_5), .POUTX(na1557_6), .POUTY1(na1557_7), .POUTY2(na1557_8),
                      .IN1(~na1530_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1530_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1529_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1544_3), .CINY1(na1556_4), .CINY2(na1556_5), .PINX(na1544_6), .PINY1(na1556_7), .PINY2(na1556_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x47y83     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1558_1 ( .COUTX(na1558_3), .COUTY1(na1558_4), .COUTY2(na1558_5), .POUTX(na1558_6), .POUTY1(na1558_7), .POUTY2(na1558_8),
                      .IN1(~na1531_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1531_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1530_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1545_3), .CINY1(na1557_4), .CINY2(na1557_5), .PINX(na1545_6), .PINY1(na1557_7), .PINY2(na1557_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x47y84     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1559_3 ( .COMP_OUT(na1559_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1559_4 ( .OUT(na1559_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1558_4), .PINX(1'b0), .PINY1(na1558_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1559_6 ( .COUTX(na1559_3), .POUTX(na1559_6), .CINX(1'b0), .CINY1(na1558_4), .CINY2(na1558_5), .PINX(1'b0), .PINY1(na1558_7),
                      .PINY2(na1558_8), .OUT1(1'b0), .OUT2(na1559_2), .COMP_OUT(na1559_3_i) );
// C_AND///AND/      x48y72     80'h00_0078_12_0000_0C88_FAAF
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1560_1 ( .OUT(na1560_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na67_1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1560_4 ( .OUT(na1560_2), .IN1(1'b1), .IN2(1'b1), .IN3(na69_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1560_6 ( .COUTY1(na1560_4), .POUTY1(na1560_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1560_1), .OUT2(na1560_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x48y73     80'h00_0018_04_2056_5888_0CCF
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1561_1 ( .OUT(na1561_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(na1548_3), .CINY1(na1560_4), .PINX(1'b0), .PINY1(na1560_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1561_3 ( .COMP_OUT(na1561_3_i), .COMB1(na1561_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1561_6 ( .COUTY1(na1561_4), .COUTY2(na1561_5), .POUTY1(na1561_7), .CINX(na1548_3), .CINY1(na1560_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1560_7), .PINY2(1'b0), .OUT1(na1561_1), .OUT2(1'b0), .COMP_OUT(na1561_3_i) );
// C_MULTFa//O_O2//      x48y74     80'h00_0018_13_A477_34A6_0CCC
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1562_1 ( .COUTX(na1562_3), .COUTY1(na1562_4), .COUTY2(na1562_5), .POUTY1(na1562_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1549_3), .CINY1(na1561_4),
                      .CINY2(na1561_5), .PINX(1'b0), .PINY1(na1561_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x48y75     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1563_1 ( .OUT(na1563_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1562_4), .PINX(1'b0), .PINY1(na1562_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1563_3 ( .COMP_OUT(na1563_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1563_4 ( .OUT(na1563_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1562_4), .PINX(1'b0), .PINY1(na1562_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1563_6 ( .COUTX(na1563_3), .COUTY1(na1563_4), .COUTY2(na1563_5), .POUTY1(na1563_7), .POUTY2(na1563_8), .CINX(1'b0), .CINY1(na1562_4),
                      .CINY2(na1562_5), .PINX(1'b0), .PINY1(na1562_7), .PINY2(1'b0), .OUT1(na1563_1), .OUT2(na1563_2), .COMP_OUT(na1563_3_i) );
// C_MULT///MULT/      x48y76     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1564_1 ( .COUTY1(na1564_4), .COUTY2(na1564_5), .POUTY1(na1564_7), .POUTY2(na1564_8), .IN1(na1523_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1523_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1522_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1551_3),
                      .CINY1(na1563_4), .CINY2(na1563_5), .PINX(na1551_6), .PINY1(na1563_7), .PINY2(na1563_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x48y77     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1565_1 ( .COUTX(na1565_3), .COUTY1(na1565_4), .COUTY2(na1565_5), .POUTX(na1565_6), .POUTY1(na1565_7), .POUTY2(na1565_8),
                      .IN1(na1524_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1524_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1523_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1552_3), .CINY1(na1564_4), .CINY2(na1564_5), .PINX(na1552_6), .PINY1(na1564_7), .PINY2(na1564_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x48y78     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1566_1 ( .COUTX(na1566_3), .COUTY1(na1566_4), .COUTY2(na1566_5), .POUTX(na1566_6), .POUTY1(na1566_7), .POUTY2(na1566_8),
                      .IN1(na1525_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1525_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1524_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1553_3), .CINY1(na1565_4), .CINY2(na1565_5), .PINX(na1553_6), .PINY1(na1565_7), .PINY2(na1565_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x48y79     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1567_1 ( .COUTX(na1567_3), .COUTY1(na1567_4), .COUTY2(na1567_5), .POUTX(na1567_6), .POUTY1(na1567_7), .POUTY2(na1567_8),
                      .IN1(na1526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1526_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1525_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1554_3), .CINY1(na1566_4), .CINY2(na1566_5), .PINX(na1554_6), .PINY1(na1566_7), .PINY2(na1566_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x48y80     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1568_1 ( .COUTX(na1568_3), .COUTY1(na1568_4), .COUTY2(na1568_5), .POUTX(na1568_6), .POUTY1(na1568_7), .POUTY2(na1568_8),
                      .IN1(na1527_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1527_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1526_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1555_3), .CINY1(na1567_4), .CINY2(na1567_5), .PINX(na1555_6), .PINY1(na1567_7), .PINY2(na1567_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x48y81     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1569_1 ( .COUTX(na1569_3), .COUTY1(na1569_4), .COUTY2(na1569_5), .POUTX(na1569_6), .POUTY1(na1569_7), .POUTY2(na1569_8),
                      .IN1(na1528_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1528_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1527_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1556_3), .CINY1(na1568_4), .CINY2(na1568_5), .PINX(na1556_6), .PINY1(na1568_7), .PINY2(na1568_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x48y82     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1570_1 ( .COUTX(na1570_3), .COUTY1(na1570_4), .COUTY2(na1570_5), .POUTX(na1570_6), .POUTY1(na1570_7), .POUTY2(na1570_8),
                      .IN1(na1529_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1529_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1528_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1557_3), .CINY1(na1569_4), .CINY2(na1569_5), .PINX(na1557_6), .PINY1(na1569_7), .PINY2(na1569_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x48y83     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1571_1 ( .COUTX(na1571_3), .COUTY1(na1571_4), .COUTY2(na1571_5), .POUTX(na1571_6), .POUTY1(na1571_7), .POUTY2(na1571_8),
                      .IN1(na1530_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1530_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1529_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1558_3), .CINY1(na1570_4), .CINY2(na1570_5), .PINX(na1558_6), .PINY1(na1570_7), .PINY2(na1570_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x48y84     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1572_1 ( .COUTX(na1572_3), .COUTY1(na1572_4), .COUTY2(na1572_5), .POUTX(na1572_6), .POUTY1(na1572_7), .POUTY2(na1572_8),
                      .IN1(na1531_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1531_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1530_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1559_3), .CINY1(na1571_4), .CINY2(na1571_5), .PINX(na1559_6), .PINY1(na1571_7), .PINY2(na1571_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x48y85     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1573_3 ( .COMP_OUT(na1573_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1573_4 ( .OUT(na1573_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1572_4), .PINX(1'b0), .PINY1(na1572_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1573_6 ( .COUTX(na1573_3), .POUTX(na1573_6), .CINX(1'b0), .CINY1(na1572_4), .CINY2(na1572_5), .PINX(1'b0), .PINY1(na1572_7),
                      .PINY2(na1572_8), .OUT1(1'b0), .OUT2(na1573_2), .COMP_OUT(na1573_3_i) );
// C_AND///AND/      x49y73     80'h00_0078_12_0000_0C88_F1F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1574_1 ( .OUT(na1574_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1051_1), .IN6(~na613_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1574_4 ( .OUT(na1574_2), .IN1(~na1051_1), .IN2(~na613_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1574_6 ( .COUTY1(na1574_4), .POUTY1(na1574_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1574_1), .OUT2(na1574_2), .COMP_OUT(1'b0) );
// C_OR//O_O1//      x49y74     80'h00_0018_04_2056_5EEE_0CC0
C_OR       #(.CPE_CFG (9'b0_0001_0110)) 
           _a1575_1 ( .OUT(na1575_1), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(na1562_3), .CINY1(na1574_4), .PINX(1'b0), .PINY1(na1574_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1575_3 ( .COMP_OUT(na1575_3_i), .COMB1(na1575_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1575_6 ( .COUTY1(na1575_4), .COUTY2(na1575_5), .POUTY1(na1575_7), .CINX(na1562_3), .CINY1(na1574_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1574_7), .PINY2(1'b0), .OUT1(na1575_1), .OUT2(1'b0), .COMP_OUT(na1575_3_i) );
// C_MULTFb//O_O2//      x49y75     80'h00_0018_13_A477_3EA6_0CCC
C_MULTFb   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1576_1 ( .COUTX(na1576_3), .COUTY1(na1576_4), .COUTY2(na1576_5), .POUTY1(na1576_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1),
                      .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1563_3), .CINY1(na1575_4),
                      .CINY2(na1575_5), .PINX(1'b0), .PINY1(na1575_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_O2/AND/      x49y76     80'h00_0078_35_A471_3C88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1577_1 ( .OUT(na1577_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1576_4), .PINX(1'b0), .PINY1(na1576_7) );
C_O_O2     #(.CPE_CFG ()) 
           _a1577_3 ( .COMP_OUT(na1577_3_i), .COMB1(1'b0), .COMB2(na1577_2) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1577_4 ( .OUT(na1577_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1576_4), .PINX(1'b0), .PINY1(na1576_7) );
C_CPlines  #(.CPE_CFG (19'h3_5A47)) 
           _a1577_6 ( .COUTX(na1577_3), .COUTY1(na1577_4), .COUTY2(na1577_5), .POUTY1(na1577_7), .POUTY2(na1577_8), .CINX(1'b0), .CINY1(na1576_4),
                      .CINY2(na1576_5), .PINX(1'b0), .PINY1(na1576_7), .PINY2(1'b0), .OUT1(na1577_1), .OUT2(na1577_2), .COMP_OUT(na1577_3_i) );
// C_MULT///MULT/      x49y77     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1578_1 ( .OUT1(na1578_1), .OUT2(na1578_2), .COUTY1(na1578_4), .COUTY2(na1578_5), .POUTY1(na1578_7), .POUTY2(na1578_8), .IN1(~na1523_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1523_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1522_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1565_3), .CINY1(na1577_4), .CINY2(na1577_5), .PINX(na1565_6), .PINY1(na1577_7), .PINY2(na1577_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x49y78     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1579_1 ( .COUTX(na1579_3), .COUTY1(na1579_4), .COUTY2(na1579_5), .POUTX(na1579_6), .POUTY1(na1579_7), .POUTY2(na1579_8),
                      .IN1(~na1524_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1524_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1523_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1566_3), .CINY1(na1578_4), .CINY2(na1578_5), .PINX(na1566_6), .PINY1(na1578_7), .PINY2(na1578_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x49y79     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1580_1 ( .COUTX(na1580_3), .COUTY1(na1580_4), .COUTY2(na1580_5), .POUTX(na1580_6), .POUTY1(na1580_7), .POUTY2(na1580_8),
                      .IN1(~na1525_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1525_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1524_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1567_3), .CINY1(na1579_4), .CINY2(na1579_5), .PINX(na1567_6), .PINY1(na1579_7), .PINY2(na1579_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x49y80     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1581_1 ( .COUTX(na1581_3), .COUTY1(na1581_4), .COUTY2(na1581_5), .POUTX(na1581_6), .POUTY1(na1581_7), .POUTY2(na1581_8),
                      .IN1(~na1526_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1526_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1525_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1568_3), .CINY1(na1580_4), .CINY2(na1580_5), .PINX(na1568_6), .PINY1(na1580_7), .PINY2(na1580_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x49y81     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1582_1 ( .COUTX(na1582_3), .COUTY1(na1582_4), .COUTY2(na1582_5), .POUTX(na1582_6), .POUTY1(na1582_7), .POUTY2(na1582_8),
                      .IN1(~na1527_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1527_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1526_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1569_3), .CINY1(na1581_4), .CINY2(na1581_5), .PINX(na1569_6), .PINY1(na1581_7), .PINY2(na1581_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x49y82     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1583_1 ( .COUTX(na1583_3), .COUTY1(na1583_4), .COUTY2(na1583_5), .POUTX(na1583_6), .POUTY1(na1583_7), .POUTY2(na1583_8),
                      .IN1(~na1528_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1528_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1527_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1570_3), .CINY1(na1582_4), .CINY2(na1582_5), .PINX(na1570_6), .PINY1(na1582_7), .PINY2(na1582_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x49y83     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1584_1 ( .COUTX(na1584_3), .COUTY1(na1584_4), .COUTY2(na1584_5), .POUTX(na1584_6), .POUTY1(na1584_7), .POUTY2(na1584_8),
                      .IN1(~na1529_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1529_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1528_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1571_3), .CINY1(na1583_4), .CINY2(na1583_5), .PINX(na1571_6), .PINY1(na1583_7), .PINY2(na1583_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x49y84     80'h00_0000_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1585_1 ( .COUTX(na1585_3), .COUTY1(na1585_4), .COUTY2(na1585_5), .POUTX(na1585_6), .POUTY1(na1585_7), .POUTY2(na1585_8),
                      .IN1(~na1530_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1530_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1529_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1572_3), .CINY1(na1584_4), .CINY2(na1584_5), .PINX(na1572_6), .PINY1(na1584_7), .PINY2(na1584_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x49y85     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1586_1 ( .COUTX(na1586_3), .COUTY1(na1586_4), .COUTY2(na1586_5), .POUTX(na1586_6), .POUTY1(na1586_7), .POUTY2(na1586_8),
                      .IN1(~na1531_2), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1531_1), .IN6(1'b1), .IN7(1'b1), .IN8(~na1530_2), .CLK(1'b0),
                      .EN(1'b0), .SR(1'b0), .CINX(na1573_3), .CINY1(na1585_4), .CINY2(na1585_5), .PINX(na1573_6), .PINY1(na1585_7), .PINY2(na1585_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x49y86     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1587_3 ( .COMP_OUT(na1587_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1587_4 ( .OUT(na1587_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1586_4), .PINX(1'b0), .PINY1(na1586_7) );
C_CPlines  #(.CPE_CFG (19'h3_9440)) 
           _a1587_6 ( .COUTX(na1587_3), .POUTX(na1587_6), .CINX(1'b0), .CINY1(na1586_4), .CINY2(na1586_5), .PINX(1'b0), .PINY1(na1586_7),
                      .PINY2(na1586_8), .OUT1(1'b0), .OUT2(na1587_2), .COMP_OUT(na1587_3_i) );
// C_AND///AND/      x50y74     80'h00_0078_12_0000_0C88_F1F1
C_AND      #(.CPE_CFG (9'b0_0000_0000)) 
           _a1588_1 ( .OUT(na1588_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(~na1051_1), .IN6(~na613_1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1588_4 ( .OUT(na1588_2), .IN1(~na1051_1), .IN2(~na613_1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h1_2000)) 
           _a1588_6 ( .COUTY1(na1588_4), .POUTY1(na1588_7), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0),
                      .OUT1(na1588_1), .OUT2(na1588_2), .COMP_OUT(1'b0) );
// C_AND//O_O1//      x50y75     80'h00_0018_04_2056_5888_0CCF
C_AND      #(.CPE_CFG (9'b0_0001_0110)) 
           _a1589_1 ( .OUT(na1589_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(na1576_3), .CINY1(na1588_4), .PINX(1'b0), .PINY1(na1588_7) );
C_O_O1     #(.CPE_CFG ()) 
           _a1589_3 ( .COMP_OUT(na1589_3_i), .COMB1(na1589_1), .COMB2(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_4205)) 
           _a1589_6 ( .COUTY1(na1589_4), .COUTY2(na1589_5), .POUTY1(na1589_7), .CINX(na1576_3), .CINY1(na1588_4), .CINY2(1'b0), .PINX(1'b0),
                      .PINY1(na1588_7), .PINY2(1'b0), .OUT1(na1589_1), .OUT2(1'b0), .COMP_OUT(na1589_3_i) );
// C_MULTFa//O_O2//      x50y76     80'h00_0018_13_A477_34A6_0CCC
C_MULTFa   #(.CPE_CFG (9'b0_0001_0111)) 
           _a1590_1 ( .COUTY1(na1590_4), .COUTY2(na1590_5), .POUTY1(na1590_7), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1),
                      .IN6(1'b1), .IN7(1'b1), .IN8(1'b1), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1577_3), .CINY1(na1589_4), .CINY2(na1589_5),
                      .PINX(1'b0), .PINY1(na1589_7), .PINY2(1'b0), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_AND//O_0/AND/      x50y77     80'h00_0078_37_A471_FC88_F0FC
C_AND      #(.CPE_CFG (9'b0_0010_0000)) 
           _a1591_1 ( .OUT(na1591_1), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b0), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1590_4), .PINX(1'b0), .PINY1(na1590_7) );
C_O_0      #(.CPE_CFG ()) 
           _a1591_3 ( .COMP_OUT(na1591_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_AND      #(.CPE_CFG (9'b0_1000_0001)) 
           _a1591_4 ( .OUT(na1591_2), .IN1(1'b1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(na1590_4), .PINX(1'b0), .PINY1(na1590_7) );
C_CPlines  #(.CPE_CFG (19'h3_7A47)) 
           _a1591_6 ( .COUTY1(na1591_4), .COUTY2(na1591_5), .POUTY1(na1591_7), .POUTY2(na1591_8), .CINX(1'b0), .CINY1(na1590_4), .CINY2(na1590_5),
                      .PINX(1'b0), .PINY1(na1590_7), .PINY2(1'b0), .OUT1(na1591_1), .OUT2(na1591_2), .COMP_OUT(na1591_3_i) );
// C_MULT///MULT/      x50y78     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1592_1 ( .OUT1(na1592_1), .OUT2(na1592_2), .COUTY1(na1592_4), .COUTY2(na1592_5), .POUTY1(na1592_7), .POUTY2(na1592_8), .IN1(na1523_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1523_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1522_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1579_3), .CINY1(na1591_4), .CINY2(na1591_5), .PINX(na1579_6), .PINY1(na1591_7), .PINY2(na1591_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x50y79     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1593_1 ( .OUT1(na1593_1), .OUT2(na1593_2), .COUTY1(na1593_4), .COUTY2(na1593_5), .POUTY1(na1593_7), .POUTY2(na1593_8), .IN1(na1524_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1524_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1523_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1580_3), .CINY1(na1592_4), .CINY2(na1592_5), .PINX(na1580_6), .PINY1(na1592_7), .PINY2(na1592_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x50y80     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1594_1 ( .OUT1(na1594_1), .OUT2(na1594_2), .COUTY1(na1594_4), .COUTY2(na1594_5), .POUTY1(na1594_7), .POUTY2(na1594_8), .IN1(na1525_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1525_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1524_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1581_3), .CINY1(na1593_4), .CINY2(na1593_5), .PINX(na1581_6), .PINY1(na1593_7), .PINY2(na1593_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x50y81     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1595_1 ( .OUT1(na1595_1), .OUT2(na1595_2), .COUTY1(na1595_4), .COUTY2(na1595_5), .POUTY1(na1595_7), .POUTY2(na1595_8), .IN1(na1526_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1526_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1525_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1582_3), .CINY1(na1594_4), .CINY2(na1594_5), .PINX(na1582_6), .PINY1(na1594_7), .PINY2(na1594_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x50y82     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1596_1 ( .OUT1(na1596_1), .OUT2(na1596_2), .COUTY1(na1596_4), .COUTY2(na1596_5), .POUTY1(na1596_7), .POUTY2(na1596_8), .IN1(na1527_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1527_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1526_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1583_3), .CINY1(na1595_4), .CINY2(na1595_5), .PINX(na1583_6), .PINY1(na1595_7), .PINY2(na1595_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x50y83     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1597_1 ( .OUT1(na1597_1), .OUT2(na1597_2), .COUTY1(na1597_4), .COUTY2(na1597_5), .POUTY1(na1597_7), .POUTY2(na1597_8), .IN1(na1528_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1528_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1527_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1584_3), .CINY1(na1596_4), .CINY2(na1596_5), .PINX(na1584_6), .PINY1(na1596_7), .PINY2(na1596_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x50y84     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1598_1 ( .OUT1(na1598_1), .OUT2(na1598_2), .COUTY1(na1598_4), .COUTY2(na1598_5), .POUTY1(na1598_7), .POUTY2(na1598_8), .IN1(na1529_2),
                      .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(na1529_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1528_2), .CLK(1'b0), .EN(1'b0),
                      .SR(1'b0), .CINX(na1585_3), .CINY1(na1597_4), .CINY2(na1597_5), .PINX(na1585_6), .PINY1(na1597_7), .PINY2(na1597_8),
                      .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x50y85     80'h00_0050_00_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0000_1100)) 
           _a1599_1 ( .COUTY1(na1599_4), .COUTY2(na1599_5), .POUTY1(na1599_7), .POUTY2(na1599_8), .IN1(na1530_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1530_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1529_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1586_3),
                      .CINY1(na1598_4), .CINY2(na1598_5), .PINX(na1586_6), .PINY1(na1598_7), .PINY2(na1598_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_MULT///MULT/      x50y86     80'h00_0010_50_003F_0C66_C8C8
C_MULT     #(.CPE_CFG (9'b0_0001_1100)) 
           _a1600_1 ( .COUTY1(na1600_4), .COUTY2(na1600_5), .POUTY1(na1600_7), .POUTY2(na1600_8), .IN1(na1531_2), .IN2(1'b1), .IN3(1'b1),
                      .IN4(1'b1), .IN5(na1531_1), .IN6(1'b1), .IN7(1'b1), .IN8(na1530_2), .CLK(1'b0), .EN(1'b0), .SR(1'b0), .CINX(na1587_3),
                      .CINY1(na1599_4), .CINY2(na1599_5), .PINX(na1587_6), .PINY1(na1599_7), .PINY2(na1599_8), .RAM_I1(1'b0), .RAM_I2(1'b0) );
// C_//O_0/OR/      x50y87     80'h00_0060_39_4401_FC0E_FF0C
C_O_0      #(.CPE_CFG ()) 
           _a1601_3 ( .COMP_OUT(na1601_3_i), .COMB1(1'b0), .COMB2(1'b0) );
C_OR       #(.CPE_CFG (9'b0_1000_0001)) 
           _a1601_4 ( .OUT(na1601_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0),
                      .CINX(1'b0), .CINY1(na1600_4), .PINX(1'b0), .PINY1(na1600_7) );
// C_///AND/      x160y25     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1602_4 ( .OUT(na1602_2), .IN1(na774_1), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1602_6 ( .RAM_O2(na1602_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1602_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y95     80'h08_0060_00_0000_0C08_FFAF
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1603_4 ( .OUT(na1603_2), .IN1(1'b1), .IN2(1'b1), .IN3(na990_1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1603_6 ( .RAM_O2(na1603_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1603_2), .COMP_OUT(1'b0) );
// C_///AND/      x1y39     80'h08_0060_00_0000_0C08_FFFA
C_AND      #(.CPE_CFG (9'b0_1000_0000)) 
           _a1604_4 ( .OUT(na1604_2), .IN1(1'b0), .IN2(1'b1), .IN3(1'b1), .IN4(1'b1), .IN5(1'b1), .IN6(1'b1), .IN7(1'b1), .IN8(1'b1),
                      .CINX(1'b0), .CINY1(1'b0), .PINX(1'b0), .PINY1(1'b0) );
C_CPlines  #(.CPE_CFG (19'h0_0000)) 
           _a1604_6 ( .RAM_O2(na1604_10), .CINX(1'b0), .CINY1(1'b0), .CINY2(1'b0), .PINX(1'b0), .PINY1(1'b0), .PINY2(1'b0), .OUT1(1'b0),
                      .OUT2(na1604_2), .COMP_OUT(1'b0) );
// C_////Bridge      x21y77     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1605_5 ( .OUT(na1605_2), .IN1(1'b0), .IN2(1'b0), .IN3(na4_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y74     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1606_5 ( .OUT(na1606_2), .IN1(1'b0), .IN2(1'b0), .IN3(na4_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y71     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1607_5 ( .OUT(na1607_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y74     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1608_5 ( .OUT(na1608_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1609_5 ( .OUT(na1609_2), .IN1(1'b0), .IN2(1'b0), .IN3(na5_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y72     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1610_5 ( .OUT(na1610_2), .IN1(na6_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1611_5 ( .OUT(na1611_2), .IN1(na6_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1612_5 ( .OUT(na1612_2), .IN1(na6_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y78     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1613_5 ( .OUT(na1613_2), .IN1(1'b0), .IN2(na7_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x27y80     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1614_5 ( .OUT(na1614_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x24y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1615_5 ( .OUT(na1615_2), .IN1(1'b0), .IN2(1'b0), .IN3(na8_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y54     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1616_5 ( .OUT(na1616_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na23_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y51     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1617_5 ( .OUT(na1617_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na23_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y47     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1618_5 ( .OUT(na1618_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na24_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y53     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1619_5 ( .OUT(na1619_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na24_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y52     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1620_5 ( .OUT(na1620_2), .IN1(1'b0), .IN2(na25_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y51     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1621_5 ( .OUT(na1621_2), .IN1(1'b0), .IN2(1'b0), .IN3(na26_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y46     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1622_5 ( .OUT(na1622_2), .IN1(1'b0), .IN2(1'b0), .IN3(na26_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y45     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1623_5 ( .OUT(na1623_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na27_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y54     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1624_5 ( .OUT(na1624_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na29_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y49     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1625_5 ( .OUT(na1625_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na31_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y56     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1626_5 ( .OUT(na1626_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na32_1), .IN8(1'b0) );
// C_////Bridge      x51y52     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1627_5 ( .OUT(na1627_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na32_2), .IN8(1'b0) );
// C_////Bridge      x40y72     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1628_5 ( .OUT(na1628_2), .IN1(na40_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y67     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1629_5 ( .OUT(na1629_2), .IN1(1'b0), .IN2(na41_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1630_5 ( .OUT(na1630_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na42_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1631_5 ( .OUT(na1631_2), .IN1(1'b0), .IN2(1'b0), .IN3(na43_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y66     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1632_5 ( .OUT(na1632_2), .IN1(na44_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1633_5 ( .OUT(na1633_2), .IN1(na45_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1634_5 ( .OUT(na1634_2), .IN1(1'b0), .IN2(1'b0), .IN3(na46_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1635_5 ( .OUT(na1635_2), .IN1(na47_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y74     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1636_5 ( .OUT(na1636_2), .IN1(1'b0), .IN2(1'b0), .IN3(na48_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y52     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1637_5 ( .OUT(na1637_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na50_1), .IN8(1'b0) );
// C_////Bridge      x56y58     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1638_5 ( .OUT(na1638_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na82_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y73     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1639_5 ( .OUT(na1639_2), .IN1(na91_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y75     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1640_5 ( .OUT(na1640_2), .IN1(1'b0), .IN2(na98_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y81     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1641_5 ( .OUT(na1641_2), .IN1(1'b0), .IN2(na98_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x22y76     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1642_5 ( .OUT(na1642_2), .IN1(1'b0), .IN2(na98_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x21y73     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1643_5 ( .OUT(na1643_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na99_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1644_5 ( .OUT(na1644_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na99_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x23y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1645_5 ( .OUT(na1645_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na99_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1646_5 ( .OUT(na1646_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na114_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1647_5 ( .OUT(na1647_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na116_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y67     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1648_5 ( .OUT(na1648_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na116_2) );
// C_////Bridge      x62y77     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1649_5 ( .OUT(na1649_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na118_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y65     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1650_5 ( .OUT(na1650_2), .IN1(1'b0), .IN2(1'b0), .IN3(na119_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y65     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1651_5 ( .OUT(na1651_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na176_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y58     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1652_5 ( .OUT(na1652_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na182_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1653_5 ( .OUT(na1653_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na184_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y64     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1654_5 ( .OUT(na1654_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na186_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y71     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1655_5 ( .OUT(na1655_2), .IN1(1'b0), .IN2(na191_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1656_5 ( .OUT(na1656_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na192_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y68     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1657_5 ( .OUT(na1657_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na195_1), .IN8(1'b0) );
// C_////Bridge      x50y67     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1658_5 ( .OUT(na1658_2), .IN1(1'b0), .IN2(na200_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y65     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1659_5 ( .OUT(na1659_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na204_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1660_5 ( .OUT(na1660_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na209_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y63     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1661_5 ( .OUT(na1661_2), .IN1(1'b0), .IN2(na213_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1662_5 ( .OUT(na1662_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na218_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y76     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1663_5 ( .OUT(na1663_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na222_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1664_5 ( .OUT(na1664_2), .IN1(1'b0), .IN2(1'b0), .IN3(na227_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y67     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1665_5 ( .OUT(na1665_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na231_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1666_5 ( .OUT(na1666_2), .IN1(na236_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x38y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1667_5 ( .OUT(na1667_2), .IN1(1'b0), .IN2(na240_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1668_5 ( .OUT(na1668_2), .IN1(na247_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y57     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1669_5 ( .OUT(na1669_2), .IN1(1'b0), .IN2(na277_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y66     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1670_5 ( .OUT(na1670_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na279_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1671_5 ( .OUT(na1671_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na292_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y70     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1672_5 ( .OUT(na1672_2), .IN1(na303_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y65     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1673_5 ( .OUT(na1673_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na329_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y64     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1674_5 ( .OUT(na1674_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na431_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y68     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1675_5 ( .OUT(na1675_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na434_2), .IN8(1'b0) );
// C_////Bridge      x39y73     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1676_5 ( .OUT(na1676_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na455_1) );
// C_////Bridge      x35y71     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1677_5 ( .OUT(na1677_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na455_2) );
// C_////Bridge      x35y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1678_5 ( .OUT(na1678_2), .IN1(1'b0), .IN2(1'b0), .IN3(na457_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y76     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1679_5 ( .OUT(na1679_2), .IN1(1'b0), .IN2(1'b0), .IN3(na457_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y71     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1680_5 ( .OUT(na1680_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na459_1) );
// C_////Bridge      x33y66     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1681_5 ( .OUT(na1681_2), .IN1(1'b0), .IN2(1'b0), .IN3(na460_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y72     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1682_5 ( .OUT(na1682_2), .IN1(1'b0), .IN2(1'b0), .IN3(na460_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x33y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1683_5 ( .OUT(na1683_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na462_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x29y63     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1684_5 ( .OUT(na1684_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na462_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y72     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1685_5 ( .OUT(na1685_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na464_1), .IN8(1'b0) );
// C_////Bridge      x41y76     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1686_5 ( .OUT(na1686_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na464_2), .IN8(1'b0) );
// C_////Bridge      x31y63     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1687_5 ( .OUT(na1687_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na466_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x35y67     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1688_5 ( .OUT(na1688_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na466_2) );
// C_////Bridge      x33y72     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1689_5 ( .OUT(na1689_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na468_1), .IN8(1'b0) );
// C_////Bridge      x35y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1690_5 ( .OUT(na1690_2), .IN1(1'b0), .IN2(1'b0), .IN3(na468_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y47     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1691_5 ( .OUT(na1691_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na583_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y50     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1692_5 ( .OUT(na1692_2), .IN1(na585_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y53     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1693_5 ( .OUT(na1693_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na590_1), .IN8(1'b0) );
// C_////Bridge      x58y55     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1694_5 ( .OUT(na1694_2), .IN1(na601_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y58     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1695_5 ( .OUT(na1695_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na603_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y53     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1696_5 ( .OUT(na1696_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na605_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y57     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1697_5 ( .OUT(na1697_2), .IN1(1'b0), .IN2(na607_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y62     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1698_5 ( .OUT(na1698_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na607_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y62     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1699_5 ( .OUT(na1699_2), .IN1(na609_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y55     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1700_5 ( .OUT(na1700_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na609_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1701_5 ( .OUT(na1701_2), .IN1(na611_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1702_5 ( .OUT(na1702_2), .IN1(na611_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y74     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1703_5 ( .OUT(na1703_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na613_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y66     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1704_5 ( .OUT(na1704_2), .IN1(na722_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y59     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1705_5 ( .OUT(na1705_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na723_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y60     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1706_5 ( .OUT(na1706_2), .IN1(na724_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y61     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1707_5 ( .OUT(na1707_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na725_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y63     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1708_5 ( .OUT(na1708_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na725_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y75     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1709_5 ( .OUT(na1709_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na726_2), .IN8(1'b0) );
// C_////Bridge      x50y72     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1710_5 ( .OUT(na1710_2), .IN1(1'b0), .IN2(na727_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y65     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1711_5 ( .OUT(na1711_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na727_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y76     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1712_5 ( .OUT(na1712_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na729_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y63     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1713_5 ( .OUT(na1713_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na729_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y75     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1714_5 ( .OUT(na1714_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na730_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y79     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1715_5 ( .OUT(na1715_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na731_1), .IN8(1'b0) );
// C_////Bridge      x61y79     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1716_5 ( .OUT(na1716_2), .IN1(1'b0), .IN2(1'b0), .IN3(na731_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1717_5 ( .OUT(na1717_2), .IN1(1'b0), .IN2(1'b0), .IN3(na731_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x41y80     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1718_5 ( .OUT(na1718_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na732_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y79     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1719_5 ( .OUT(na1719_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na733_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y69     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1720_5 ( .OUT(na1720_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na733_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1721_5 ( .OUT(na1721_2), .IN1(na734_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1722_5 ( .OUT(na1722_2), .IN1(na734_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y82     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1723_5 ( .OUT(na1723_2), .IN1(na734_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y47     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1724_5 ( .OUT(na1724_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na775_1) );
// C_////Bridge      x55y49     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1725_5 ( .OUT(na1725_2), .IN1(1'b0), .IN2(1'b0), .IN3(na777_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y49     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1726_5 ( .OUT(na1726_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na779_1) );
// C_////Bridge      x49y49     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1727_5 ( .OUT(na1727_2), .IN1(1'b0), .IN2(1'b0), .IN3(na781_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y51     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1728_5 ( .OUT(na1728_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na783_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y51     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1729_5 ( .OUT(na1729_2), .IN1(1'b0), .IN2(1'b0), .IN3(na785_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y53     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1730_5 ( .OUT(na1730_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na787_1) );
// C_////Bridge      x55y53     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1731_5 ( .OUT(na1731_2), .IN1(1'b0), .IN2(1'b0), .IN3(na789_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x53y55     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1732_5 ( .OUT(na1732_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na791_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y55     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1733_5 ( .OUT(na1733_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na793_1), .IN8(1'b0) );
// C_////Bridge      x53y61     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1734_5 ( .OUT(na1734_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na795_1) );
// C_////Bridge      x55y57     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1735_5 ( .OUT(na1735_2), .IN1(1'b0), .IN2(1'b0), .IN3(na797_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y63     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1736_5 ( .OUT(na1736_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na799_1) );
// C_////Bridge      x53y59     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1737_5 ( .OUT(na1737_2), .IN1(1'b0), .IN2(1'b0), .IN3(na801_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x25y70     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1738_5 ( .OUT(na1738_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na862_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y47     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1739_5 ( .OUT(na1739_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na866_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y50     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1740_5 ( .OUT(na1740_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na866_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y45     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1741_5 ( .OUT(na1741_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na866_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x51y46     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1742_5 ( .OUT(na1742_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na868_1), .IN8(1'b0) );
// C_////Bridge      x30y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1743_5 ( .OUT(na1743_2), .IN1(1'b0), .IN2(na871_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x28y76     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1744_5 ( .OUT(na1744_2), .IN1(1'b0), .IN2(na871_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x31y75     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1745_5 ( .OUT(na1745_2), .IN1(1'b0), .IN2(na871_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x32y78     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1746_5 ( .OUT(na1746_2), .IN1(1'b0), .IN2(na871_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x61y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1747_5 ( .OUT(na1747_2), .IN1(1'b0), .IN2(na889_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y70     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1748_5 ( .OUT(na1748_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na891_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y69     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1749_5 ( .OUT(na1749_2), .IN1(na895_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1750_5 ( .OUT(na1750_2), .IN1(na895_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y70     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1751_5 ( .OUT(na1751_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na895_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y74     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1752_5 ( .OUT(na1752_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na897_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y78     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1753_5 ( .OUT(na1753_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na897_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y75     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1754_5 ( .OUT(na1754_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na899_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y77     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1755_5 ( .OUT(na1755_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na899_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y73     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1756_5 ( .OUT(na1756_2), .IN1(1'b0), .IN2(na901_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y79     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1757_5 ( .OUT(na1757_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na901_2), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y76     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1758_5 ( .OUT(na1758_2), .IN1(na931_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x49y71     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1759_5 ( .OUT(na1759_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na933_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x44y75     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1760_5 ( .OUT(na1760_2), .IN1(1'b0), .IN2(na935_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x42y80     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1761_5 ( .OUT(na1761_2), .IN1(na937_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y59     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1762_5 ( .OUT(na1762_2), .IN1(1'b0), .IN2(na942_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y64     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1763_5 ( .OUT(na1763_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na944_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y57     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1764_5 ( .OUT(na1764_2), .IN1(1'b0), .IN2(na946_2), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y65     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1765_5 ( .OUT(na1765_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na949_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x48y47     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1766_5 ( .OUT(na1766_2), .IN1(na951_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y63     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1767_5 ( .OUT(na1767_2), .IN1(1'b0), .IN2(na953_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x46y62     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1768_5 ( .OUT(na1768_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na955_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y73     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1769_5 ( .OUT(na1769_2), .IN1(1'b0), .IN2(1'b0), .IN3(na958_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1770_5 ( .OUT(na1770_2), .IN1(1'b0), .IN2(1'b0), .IN3(na958_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y77     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1771_5 ( .OUT(na1771_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na960_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y76     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1772_5 ( .OUT(na1772_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na960_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y81     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1773_5 ( .OUT(na1773_2), .IN1(1'b0), .IN2(1'b0), .IN3(na962_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1774_5 ( .OUT(na1774_2), .IN1(1'b0), .IN2(1'b0), .IN3(na962_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y80     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1775_5 ( .OUT(na1775_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na963_1) );
// C_////Bridge      x57y68     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1776_5 ( .OUT(na1776_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na965_1), .IN8(1'b0) );
// C_////Bridge      x57y67     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1777_5 ( .OUT(na1777_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na967_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y70     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1778_5 ( .OUT(na1778_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na967_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y72     80'h00_00A6_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1779_5 ( .OUT(na1779_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(na969_1), .IN8(1'b0) );
// C_////Bridge      x63y75     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1780_5 ( .OUT(na1780_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na971_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y74     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1781_5 ( .OUT(na1781_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na971_1), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x57y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1782_5 ( .OUT(na1782_2), .IN1(na974_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1783_5 ( .OUT(na1783_2), .IN1(na974_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y78     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1784_5 ( .OUT(na1784_2), .IN1(na974_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x59y71     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1785_5 ( .OUT(na1785_2), .IN1(1'b0), .IN2(na976_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y67     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1786_5 ( .OUT(na1786_2), .IN1(1'b0), .IN2(na976_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y80     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1787_5 ( .OUT(na1787_2), .IN1(1'b0), .IN2(na976_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y78     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1788_5 ( .OUT(na1788_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na978_1), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y76     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1789_5 ( .OUT(na1789_2), .IN1(1'b0), .IN2(na979_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y79     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1790_5 ( .OUT(na1790_2), .IN1(1'b0), .IN2(na979_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y74     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1791_5 ( .OUT(na1791_2), .IN1(1'b0), .IN2(na979_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1792_5 ( .OUT(na1792_2), .IN1(1'b0), .IN2(na983_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y69     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1793_5 ( .OUT(na1793_2), .IN1(1'b0), .IN2(na983_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y67     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1794_5 ( .OUT(na1794_2), .IN1(na985_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x62y72     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1795_5 ( .OUT(na1795_2), .IN1(na985_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y68     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1796_5 ( .OUT(na1796_2), .IN1(1'b0), .IN2(na987_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x60y71     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1797_5 ( .OUT(na1797_2), .IN1(1'b0), .IN2(na987_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x58y64     80'h00_00A1_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1798_5 ( .OUT(na1798_2), .IN1(1'b0), .IN2(na987_1), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x26y77     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1799_5 ( .OUT(na1799_2), .IN1(na1041_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x34y78     80'h00_00A4_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1800_5 ( .OUT(na1800_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(na1055_2), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y68     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1801_5 ( .OUT(na1801_2), .IN1(na1075_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x47y65     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1802_5 ( .OUT(na1802_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1076_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x40y73     80'h00_00A5_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1803_5 ( .OUT(na1803_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(na1087_1), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x36y74     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1804_5 ( .OUT(na1804_2), .IN1(na1090_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x50y58     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1805_5 ( .OUT(na1805_2), .IN1(na1095_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x55y75     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1806_5 ( .OUT(na1806_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1112_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x52y75     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1807_5 ( .OUT(na1807_2), .IN1(na1114_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x56y73     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1808_5 ( .OUT(na1808_2), .IN1(na1128_1), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x54y64     80'h00_00A0_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1809_5 ( .OUT(na1809_2), .IN1(na1578_2), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x39y75     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1810_5 ( .OUT(na1810_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1592_1) );
// C_////Bridge      x33y69     80'h00_00A7_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1811_5 ( .OUT(na1811_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(na1592_2) );
// C_////Bridge      x39y78     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1812_5 ( .OUT(na1812_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1593_1), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x45y70     80'h00_00A2_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1813_5 ( .OUT(na1813_2), .IN1(1'b0), .IN2(1'b0), .IN3(na1593_2), .IN4(1'b0), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
// C_////Bridge      x37y78     80'h00_00A3_00_0000_0C00_FFFF
C_Bridge   #(.CPE_CFG (9'bX_0000_1001)) 
           _a1814_5 ( .OUT(na1814_2), .IN1(1'b0), .IN2(1'b0), .IN3(1'b0), .IN4(na1598_2), .IN5(1'b0), .IN6(1'b0), .IN7(1'b0), .IN8(1'b0) );
endmodule
